module CHIP_TOP(
    
    input       sys_clk             ,
    input       sys_rst_n           ,

    output      led_test            

);
//=================================================================================
// Parameter declaration
//=================================================================================


//=================================================================================
// Signal declaration
//=================================================================================


//=================================================================================
// Body
//=================================================================================

riscv_core      u_riscv_core(
    //system signal
    .sys_clk        ( sys_clk       ),
    .sys_rst_n      ( sys_rst_n     ),
    .led_test       ( led_test      )
);

endmodule
