/*
     Copyright (c) 2023 SMIC             
     Filename:      S55NLLGSPH_X512Y16D32.lef
     IP code:       S55NLLGSPH
     Version:       1.1.a
     CreateDate:    2023-2-15        
                    
    LEF for General Single-PORT SRAM
    SMIC 55nm LL Logic Process

    Configuration: -instname S55NLLGSPH_X512Y16D32 -rows 512 -bits 32 -mux 16 
    Redundancy: Off
    Bit-Write: Off
*/

# DISCLAIMER                                                                      
#                                                                                   
#   SMIC hereby provides the quality information to you but makes no claims,      
# promises or guarantees about the accuracy, completeness, or adequacy of the     
# information herein. The information contained herein is provided on an "AS IS"  
# basis without any warranty, and SMIC assumes no obligation to provide support   
# of any kind or otherwise maintain the information.                                
#   SMIC disclaims any representation that the information does not infringe any  
# intellectual property rights or proprietary rights of any third parties. SMIC   
# makes no other warranty, whether express, implied or statutory as to any        
# matter whatsoever, including but not limited to the accuracy or sufficiency of  
# any information or the merchantability and fitness for a particular purpose.    
# Neither SMIC nor any of its representatives shall be liable for any cause of    
# action incurred to connect to this service.                                       
#                                                                                 
# STATEMENT OF USE AND CONFIDENTIALITY                                              
#                                                                                   
#   The following/attached material contains confidential and proprietary           
# information of SMIC. This material is based upon information which SMIC           
# considers reliable, but SMIC neither represents nor warrants that such          
# information is accurate or complete, and it must not be relied upon as such.    
# This information was prepared for informational purposes and is for the use     
# by SMIC's customer only. SMIC reserves the right to make changes in the           
# information at any time without notice.                                           
#   No part of this information may be reproduced, transmitted, transcribed,        
# stored in a retrieval system, or translated into any human or computer           
# language, in any form or by any means, electronic, mechanical, magnetic,          
# optical, chemical, manual, or otherwise, without the prior written consent of   
# SMIC. Any unauthorized use or disclosure of this material is strictly             
# prohibited and may be unlawful. By accepting this material, the receiving         
# party shall be deemed to have acknowledged, accepted, and agreed to be bound    
# by the foregoing limitations and restrictions. Thank you.                         
#                                                                                   

VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO S55NLLGSPH_X512Y16D32
 CLASS BLOCK ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SIZE 569.26 BY 307.045 ;

 PIN A[11]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 270.025 0 270.225 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 270.025 0 270.225 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 270.025 0 270.225 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END A[11]

 PIN A[12]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 270.425 0 270.625 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 270.425 0 270.625 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 270.425 0 270.625 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END A[12]

 PIN A[9]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 270.825 0 271.025 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 270.825 0 271.025 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 270.825 0 271.025 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END A[9]

 PIN A[10]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 271.225 0 271.425 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 271.225 0 271.425 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 271.225 0 271.425 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END A[10]

 PIN A[3]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 276.905 0 277.105 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 276.905 0 277.105 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 276.905 0 277.105 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END A[3]

 PIN A[7]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 277.305 0 277.505 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 277.305 0 277.505 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 277.305 0 277.505 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END A[7]

 PIN A[8]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 280.205 0 280.405 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 280.205 0 280.405 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 280.205 0 280.405 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END A[8]

 PIN A[4]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 280.655 0 280.855 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 280.655 0 280.855 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 280.655 0 280.855 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END A[4]

 PIN A[6]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 281.105 0 281.305 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 281.105 0 281.305 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 281.105 0 281.305 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END A[6]

 PIN CEN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 281.555 0 281.755 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 281.555 0 281.755 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 281.555 0 281.755 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END CEN

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 282.01 0 282.21 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 282.01 0 282.21 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 282.01 0 282.21 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END CLK

 PIN A[5]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 288.395 0 288.595 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 288.395 0 288.595 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 288.395 0 288.595 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END A[5]

 PIN A[0]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 288.795 0 288.995 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 288.795 0 288.995 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 288.795 0 288.995 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END A[0]

 PIN A[1]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 289.195 0 289.395 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 289.195 0 289.395 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 289.195 0 289.395 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END A[1]

 PIN WEN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 292.18 0 292.38 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 292.18 0 292.38 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 292.18 0 292.38 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END WEN

 PIN A[2]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 298.195 0 298.395 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 298.195 0 298.395 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 298.195 0 298.395 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END A[2]

 PIN Q[0]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 9.155 0 9.355 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 9.155 0 9.355 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 9.155 0 9.355 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[0]

 PIN D[0]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 9.755 0 9.955 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 9.755 0 9.955 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 9.755 0 9.955 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[0]

 PIN D[1]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 25.955 0 26.155 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 25.955 0 26.155 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 25.955 0 26.155 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[1]

 PIN Q[1]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 26.555 0 26.755 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 26.555 0 26.755 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 26.555 0 26.755 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[1]

 PIN Q[2]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 42.755 0 42.955 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 42.755 0 42.955 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 42.755 0 42.955 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[2]

 PIN D[2]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 43.355 0 43.555 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 43.355 0 43.555 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 43.355 0 43.555 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[2]

 PIN D[3]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 59.555 0 59.755 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 59.555 0 59.755 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 59.555 0 59.755 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[3]

 PIN Q[3]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 60.155 0 60.355 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 60.155 0 60.355 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 60.155 0 60.355 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[3]

 PIN Q[4]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 76.355 0 76.555 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 76.355 0 76.555 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 76.355 0 76.555 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[4]

 PIN D[4]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 76.955 0 77.155 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 76.955 0 77.155 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 76.955 0 77.155 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[4]

 PIN D[5]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 93.155 0 93.355 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 93.155 0 93.355 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 93.155 0 93.355 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[5]

 PIN Q[5]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 93.755 0 93.955 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 93.755 0 93.955 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 93.755 0 93.955 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[5]

 PIN Q[6]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 109.955 0 110.155 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 109.955 0 110.155 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 109.955 0 110.155 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[6]

 PIN D[6]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 110.555 0 110.755 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 110.555 0 110.755 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 110.555 0 110.755 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[6]

 PIN D[7]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 126.755 0 126.955 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 126.755 0 126.955 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 126.755 0 126.955 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[7]

 PIN Q[7]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 127.355 0 127.555 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 127.355 0 127.555 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 127.355 0 127.555 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[7]

 PIN Q[8]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 143.555 0 143.755 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 143.555 0 143.755 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 143.555 0 143.755 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[8]

 PIN D[8]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 144.155 0 144.355 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 144.155 0 144.355 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 144.155 0 144.355 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[8]

 PIN D[9]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 160.355 0 160.555 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 160.355 0 160.555 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 160.355 0 160.555 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[9]

 PIN Q[9]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 160.955 0 161.155 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 160.955 0 161.155 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 160.955 0 161.155 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[9]

 PIN Q[10]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 177.155 0 177.355 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 177.155 0 177.355 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 177.155 0 177.355 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[10]

 PIN D[10]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 177.755 0 177.955 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 177.755 0 177.955 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 177.755 0 177.955 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[10]

 PIN D[11]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 193.955 0 194.155 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 193.955 0 194.155 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 193.955 0 194.155 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[11]

 PIN Q[11]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 194.555 0 194.755 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 194.555 0 194.755 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 194.555 0 194.755 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[11]

 PIN Q[12]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 210.755 0 210.955 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 210.755 0 210.955 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 210.755 0 210.955 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[12]

 PIN D[12]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 211.355 0 211.555 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 211.355 0 211.555 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 211.355 0 211.555 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[12]

 PIN D[13]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 227.555 0 227.755 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 227.555 0 227.755 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 227.555 0 227.755 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[13]

 PIN Q[13]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 228.155 0 228.355 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 228.155 0 228.355 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 228.155 0 228.355 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[13]

 PIN Q[14]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 244.355 0 244.555 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 244.355 0 244.555 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 244.355 0 244.555 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[14]

 PIN D[14]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 244.955 0 245.155 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 244.955 0 245.155 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 244.955 0 245.155 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[14]

 PIN D[15]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 261.155 0 261.355 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 261.155 0 261.355 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 261.155 0 261.355 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[15]

 PIN Q[15]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 261.755 0 261.955 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 261.755 0 261.955 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 261.755 0 261.955 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[15]

 PIN Q[16]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 307.305 0 307.505 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 307.305 0 307.505 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 307.305 0 307.505 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[16]

 PIN D[16]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 307.905 0 308.105 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 307.905 0 308.105 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 307.905 0 308.105 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[16]

 PIN D[17]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 324.105 0 324.305 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 324.105 0 324.305 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 324.105 0 324.305 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[17]

 PIN Q[17]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 324.705 0 324.905 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 324.705 0 324.905 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 324.705 0 324.905 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[17]

 PIN Q[18]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 340.905 0 341.105 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 340.905 0 341.105 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 340.905 0 341.105 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[18]

 PIN D[18]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 341.505 0 341.705 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 341.505 0 341.705 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 341.505 0 341.705 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[18]

 PIN D[19]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 357.705 0 357.905 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 357.705 0 357.905 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 357.705 0 357.905 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[19]

 PIN Q[19]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 358.305 0 358.505 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 358.305 0 358.505 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 358.305 0 358.505 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[19]

 PIN Q[20]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 374.505 0 374.705 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 374.505 0 374.705 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 374.505 0 374.705 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[20]

 PIN D[20]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 375.105 0 375.305 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 375.105 0 375.305 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 375.105 0 375.305 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[20]

 PIN D[21]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 391.305 0 391.505 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 391.305 0 391.505 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 391.305 0 391.505 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[21]

 PIN Q[21]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 391.905 0 392.105 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 391.905 0 392.105 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 391.905 0 392.105 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[21]

 PIN Q[22]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 408.105 0 408.305 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 408.105 0 408.305 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 408.105 0 408.305 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[22]

 PIN D[22]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 408.705 0 408.905 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 408.705 0 408.905 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 408.705 0 408.905 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[22]

 PIN D[23]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 424.905 0 425.105 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 424.905 0 425.105 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 424.905 0 425.105 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[23]

 PIN Q[23]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 425.505 0 425.705 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 425.505 0 425.705 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 425.505 0 425.705 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[23]

 PIN Q[24]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 441.705 0 441.905 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 441.705 0 441.905 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 441.705 0 441.905 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[24]

 PIN D[24]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 442.305 0 442.505 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 442.305 0 442.505 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 442.305 0 442.505 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[24]

 PIN D[25]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 458.505 0 458.705 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 458.505 0 458.705 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 458.505 0 458.705 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[25]

 PIN Q[25]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 459.105 0 459.305 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 459.105 0 459.305 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 459.105 0 459.305 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[25]

 PIN Q[26]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 475.305 0 475.505 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 475.305 0 475.505 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 475.305 0 475.505 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[26]

 PIN D[26]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 475.905 0 476.105 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 475.905 0 476.105 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 475.905 0 476.105 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[26]

 PIN D[27]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 492.105 0 492.305 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 492.105 0 492.305 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 492.105 0 492.305 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[27]

 PIN Q[27]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 492.705 0 492.905 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 492.705 0 492.905 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 492.705 0 492.905 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[27]

 PIN Q[28]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 508.905 0 509.105 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 508.905 0 509.105 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 508.905 0 509.105 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[28]

 PIN D[28]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 509.505 0 509.705 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 509.505 0 509.705 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 509.505 0 509.705 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[28]

 PIN D[29]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 525.705 0 525.905 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 525.705 0 525.905 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 525.705 0 525.905 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[29]

 PIN Q[29]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 526.305 0 526.505 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 526.305 0 526.505 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 526.305 0 526.505 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[29]

 PIN Q[30]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 542.505 0 542.705 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 542.505 0 542.705 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 542.505 0 542.705 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[30]

 PIN D[30]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 543.105 0 543.305 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 543.105 0 543.305 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 543.105 0 543.305 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[30]

 PIN D[31]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 559.305 0 559.505 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 559.305 0 559.505 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 559.305 0 559.505 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END D[31]

 PIN Q[31]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 559.905 0 560.105 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 559.905 0 560.105 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 559.905 0 560.105 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END Q[31]


 PIN VDD
 USE POWER ;
 PORT
 LAYER M4 ;
 RECT 2.105 0 4.305 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 10.505 0 12.705 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 23.205 0 25.405 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 31.605 0 33.805 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 35.705 0 37.905 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 44.105 0 46.305 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 56.805 0 59.005 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 65.205 0 67.405 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 69.305 0 71.505 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 77.705 0 79.905 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 90.405 0 92.605 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 98.805 0 101.005 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 102.905 0 105.105 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 111.305 0 113.505 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 124.005 0 126.205 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 132.405 0 134.605 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 136.505 0 138.705 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 144.905 0 147.105 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 157.605 0 159.805 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 166.005 0 168.205 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 170.105 0 172.305 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 178.505 0 180.705 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 191.205 0 193.405 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 199.605 0 201.805 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 203.705 0 205.905 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 212.105 0 214.305 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 224.805 0 227.005 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 233.205 0 235.405 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 237.305 0 239.505 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 245.705 0 247.905 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 258.405 0 260.605 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 266.805 0 269.005 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 272.305 0 274.205 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 277.905 0 279.805 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 285.995 0 287.995 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 289.795 0 291.795 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 295.18 0 297.18 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 300.255 0 302.455 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 308.655 0 310.855 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 321.355 0 323.555 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 329.755 0 331.955 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 333.855 0 336.055 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 342.255 0 344.455 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 354.955 0 357.155 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 363.355 0 365.555 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 367.455 0 369.655 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 375.855 0 378.055 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 388.555 0 390.755 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 396.955 0 399.155 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 401.055 0 403.255 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 409.455 0 411.655 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 422.155 0 424.355 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 430.555 0 432.755 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 434.655 0 436.855 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 443.055 0 445.255 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 455.755 0 457.955 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 464.155 0 466.355 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 468.255 0 470.455 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 476.655 0 478.855 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 489.355 0 491.555 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 497.755 0 499.955 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 501.855 0 504.055 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 510.255 0 512.455 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 522.955 0 525.155 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 531.355 0 533.555 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 535.455 0 537.655 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 543.855 0 546.055 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 556.555 0 558.755 307.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 564.955 0 567.155 307.045 ;    
 END 
 END VDD

 PIN VSS
 USE GROUND ;
 PORT
 LAYER M4 ;
 RECT 6.405 0 8.605 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 14.805 0 17.005 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 18.905 0 21.105 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 27.305 0 29.505 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 40.005 0 42.205 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 48.405 0 50.605 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 52.505 0 54.705 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 60.905 0 63.105 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 73.605 0 75.805 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 82.005 0 84.205 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 86.105 0 88.305 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 94.505 0 96.705 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 107.205 0 109.405 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 115.605 0 117.805 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 119.705 0 121.905 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 128.105 0 130.305 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 140.805 0 143.005 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 149.205 0 151.405 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 153.305 0 155.505 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 161.705 0 163.905 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 174.405 0 176.605 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 182.805 0 185.005 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 186.905 0 189.105 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 195.305 0 197.505 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 208.005 0 210.205 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 216.405 0 218.605 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 220.505 0 222.705 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 228.905 0 231.105 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 241.605 0 243.805 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 250.005 0 252.205 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 254.105 0 256.305 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 262.505 0 264.705 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 274.605 0 276.505 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 283.595 0 285.595 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 292.78 0 294.78 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 304.555 0 306.755 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 312.955 0 315.155 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 317.055 0 319.255 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 325.455 0 327.655 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 338.155 0 340.355 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 346.555 0 348.755 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 350.655 0 352.855 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 359.055 0 361.255 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 371.755 0 373.955 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 380.155 0 382.355 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 384.255 0 386.455 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 392.655 0 394.855 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 405.355 0 407.555 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 413.755 0 415.955 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 417.855 0 420.055 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 426.255 0 428.455 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 438.955 0 441.155 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 447.355 0 449.555 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 451.455 0 453.655 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 459.855 0 462.055 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 472.555 0 474.755 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 480.955 0 483.155 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 485.055 0 487.255 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 493.455 0 495.655 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 506.155 0 508.355 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 514.555 0 516.755 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 518.655 0 520.855 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 527.055 0 529.255 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 539.755 0 541.955 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 548.155 0 550.355 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 552.255 0 554.455 307.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 560.655 0 562.855 307.045 ;      
 END
 END VSS

 OBS
 LAYER M1 ;
 RECT 0 0 9.065 0.57 ;
 RECT 9.445 0 9.665 0.57 ;
 RECT 10.045 0 25.865 0.57 ;
 RECT 26.245 0 26.465 0.57 ;
 RECT 26.845 0 42.665 0.57 ;
 RECT 43.045 0 43.265 0.57 ;
 RECT 43.645 0 59.465 0.57 ;
 RECT 59.845 0 60.065 0.57 ;
 RECT 60.445 0 76.265 0.57 ;
 RECT 76.645 0 76.865 0.57 ;
 RECT 77.245 0 93.065 0.57 ;
 RECT 93.445 0 93.665 0.57 ;
 RECT 94.045 0 109.865 0.57 ;
 RECT 110.245 0 110.465 0.57 ;
 RECT 110.845 0 126.665 0.57 ;
 RECT 127.045 0 127.265 0.57 ;
 RECT 127.645 0 143.465 0.57 ;
 RECT 143.845 0 144.065 0.57 ;
 RECT 144.445 0 160.265 0.57 ;
 RECT 160.645 0 160.865 0.57 ;
 RECT 161.245 0 177.065 0.57 ;
 RECT 177.445 0 177.665 0.57 ;
 RECT 178.045 0 193.865 0.57 ;
 RECT 194.245 0 194.465 0.57 ;
 RECT 194.845 0 210.665 0.57 ;
 RECT 211.045 0 211.265 0.57 ;
 RECT 211.645 0 227.465 0.57 ;
 RECT 227.845 0 228.065 0.57 ;
 RECT 228.445 0 244.265 0.57 ;
 RECT 244.645 0 244.865 0.57 ;
 RECT 245.245 0 261.065 0.57 ;
 RECT 261.445 0 261.665 0.57 ;
 RECT 262.045 0 269.935 0.57 ;
 RECT 271.515 0 276.815 0.57 ;
 RECT 277.595 0 280.115 0.57 ;
 RECT 282.3 0 288.305 0.57 ;
 RECT 289.485 0 292.09 0.57 ;
 RECT 292.47 0 298.105 0.57 ;
 RECT 298.485 0 307.215 0.57 ;
 RECT 307.595 0 307.815 0.57 ;
 RECT 308.195 0 324.015 0.57 ;
 RECT 324.395 0 324.615 0.57 ;
 RECT 324.995 0 340.815 0.57 ;
 RECT 341.195 0 341.415 0.57 ;
 RECT 341.795 0 357.615 0.57 ;
 RECT 357.995 0 358.215 0.57 ;
 RECT 358.595 0 374.415 0.57 ;
 RECT 374.795 0 375.015 0.57 ;
 RECT 375.395 0 391.215 0.57 ;
 RECT 391.595 0 391.815 0.57 ;
 RECT 392.195 0 408.015 0.57 ;
 RECT 408.395 0 408.615 0.57 ;
 RECT 408.995 0 424.815 0.57 ;
 RECT 425.195 0 425.415 0.57 ;
 RECT 425.795 0 441.615 0.57 ;
 RECT 441.995 0 442.215 0.57 ;
 RECT 442.595 0 458.415 0.57 ;
 RECT 458.795 0 459.015 0.57 ;
 RECT 459.395 0 475.215 0.57 ;
 RECT 475.595 0 475.815 0.57 ;
 RECT 476.195 0 492.015 0.57 ;
 RECT 492.395 0 492.615 0.57 ;
 RECT 492.995 0 508.815 0.57 ;
 RECT 509.195 0 509.415 0.57 ;
 RECT 509.795 0 525.615 0.57 ;
 RECT 525.995 0 526.215 0.57 ;
 RECT 526.595 0 542.415 0.57 ;
 RECT 542.795 0 543.015 0.57 ;
 RECT 543.395 0 559.215 0.57 ;
 RECT 559.595 0 559.815 0.57 ;
 RECT 560.195 0 569.26 0.57 ;
 RECT 0 0.57 569.26 307.045 ;
 LAYER M2 ;
 RECT 0 0 9.055 0.58 ;
 RECT 9.455 0 9.655 0.58 ;
 RECT 10.055 0 25.855 0.58 ;
 RECT 26.255 0 26.455 0.58 ;
 RECT 26.855 0 42.655 0.58 ;
 RECT 43.055 0 43.255 0.58 ;
 RECT 43.655 0 59.455 0.58 ;
 RECT 59.855 0 60.055 0.58 ;
 RECT 60.455 0 76.255 0.58 ;
 RECT 76.655 0 76.855 0.58 ;
 RECT 77.255 0 93.055 0.58 ;
 RECT 93.455 0 93.655 0.58 ;
 RECT 94.055 0 109.855 0.58 ;
 RECT 110.255 0 110.455 0.58 ;
 RECT 110.855 0 126.655 0.58 ;
 RECT 127.055 0 127.255 0.58 ;
 RECT 127.655 0 143.455 0.58 ;
 RECT 143.855 0 144.055 0.58 ;
 RECT 144.455 0 160.255 0.58 ;
 RECT 160.655 0 160.855 0.58 ;
 RECT 161.255 0 177.055 0.58 ;
 RECT 177.455 0 177.655 0.58 ;
 RECT 178.055 0 193.855 0.58 ;
 RECT 194.255 0 194.455 0.58 ;
 RECT 194.855 0 210.655 0.58 ;
 RECT 211.055 0 211.255 0.58 ;
 RECT 211.655 0 227.455 0.58 ;
 RECT 227.855 0 228.055 0.58 ;
 RECT 228.455 0 244.255 0.58 ;
 RECT 244.655 0 244.855 0.58 ;
 RECT 245.255 0 261.055 0.58 ;
 RECT 261.455 0 261.655 0.58 ;
 RECT 262.055 0 269.925 0.58 ;
 RECT 271.525 0 276.805 0.58 ;
 RECT 277.605 0 280.105 0.58 ;
 RECT 282.31 0 288.295 0.58 ;
 RECT 289.495 0 292.08 0.58 ;
 RECT 292.48 0 298.095 0.58 ;
 RECT 298.495 0 307.205 0.58 ;
 RECT 307.605 0 307.805 0.58 ;
 RECT 308.205 0 324.005 0.58 ;
 RECT 324.405 0 324.605 0.58 ;
 RECT 325.005 0 340.805 0.58 ;
 RECT 341.205 0 341.405 0.58 ;
 RECT 341.805 0 357.605 0.58 ;
 RECT 358.005 0 358.205 0.58 ;
 RECT 358.605 0 374.405 0.58 ;
 RECT 374.805 0 375.005 0.58 ;
 RECT 375.405 0 391.205 0.58 ;
 RECT 391.605 0 391.805 0.58 ;
 RECT 392.205 0 408.005 0.58 ;
 RECT 408.405 0 408.605 0.58 ;
 RECT 409.005 0 424.805 0.58 ;
 RECT 425.205 0 425.405 0.58 ;
 RECT 425.805 0 441.605 0.58 ;
 RECT 442.005 0 442.205 0.58 ;
 RECT 442.605 0 458.405 0.58 ;
 RECT 458.805 0 459.005 0.58 ;
 RECT 459.405 0 475.205 0.58 ;
 RECT 475.605 0 475.805 0.58 ;
 RECT 476.205 0 492.005 0.58 ;
 RECT 492.405 0 492.605 0.58 ;
 RECT 493.005 0 508.805 0.58 ;
 RECT 509.205 0 509.405 0.58 ;
 RECT 509.805 0 525.605 0.58 ;
 RECT 526.005 0 526.205 0.58 ;
 RECT 526.605 0 542.405 0.58 ;
 RECT 542.805 0 543.005 0.58 ;
 RECT 543.405 0 559.205 0.58 ;
 RECT 559.605 0 559.805 0.58 ;
 RECT 560.205 0 569.26 0.58 ;
 RECT 0 0.58 569.26 307.045 ;
 LAYER M3 ;
 RECT 0 0 9.055 0.58 ;
 RECT 9.455 0 9.655 0.58 ;
 RECT 10.055 0 25.855 0.58 ;
 RECT 26.255 0 26.455 0.58 ;
 RECT 26.855 0 42.655 0.58 ;
 RECT 43.055 0 43.255 0.58 ;
 RECT 43.655 0 59.455 0.58 ;
 RECT 59.855 0 60.055 0.58 ;
 RECT 60.455 0 76.255 0.58 ;
 RECT 76.655 0 76.855 0.58 ;
 RECT 77.255 0 93.055 0.58 ;
 RECT 93.455 0 93.655 0.58 ;
 RECT 94.055 0 109.855 0.58 ;
 RECT 110.255 0 110.455 0.58 ;
 RECT 110.855 0 126.655 0.58 ;
 RECT 127.055 0 127.255 0.58 ;
 RECT 127.655 0 143.455 0.58 ;
 RECT 143.855 0 144.055 0.58 ;
 RECT 144.455 0 160.255 0.58 ;
 RECT 160.655 0 160.855 0.58 ;
 RECT 161.255 0 177.055 0.58 ;
 RECT 177.455 0 177.655 0.58 ;
 RECT 178.055 0 193.855 0.58 ;
 RECT 194.255 0 194.455 0.58 ;
 RECT 194.855 0 210.655 0.58 ;
 RECT 211.055 0 211.255 0.58 ;
 RECT 211.655 0 227.455 0.58 ;
 RECT 227.855 0 228.055 0.58 ;
 RECT 228.455 0 244.255 0.58 ;
 RECT 244.655 0 244.855 0.58 ;
 RECT 245.255 0 261.055 0.58 ;
 RECT 261.455 0 261.655 0.58 ;
 RECT 262.055 0 269.925 0.58 ;
 RECT 271.525 0 276.805 0.58 ;
 RECT 277.605 0 280.105 0.58 ;
 RECT 282.31 0 288.295 0.58 ;
 RECT 289.495 0 292.08 0.58 ;
 RECT 292.48 0 298.095 0.58 ;
 RECT 298.495 0 307.205 0.58 ;
 RECT 307.605 0 307.805 0.58 ;
 RECT 308.205 0 324.005 0.58 ;
 RECT 324.405 0 324.605 0.58 ;
 RECT 325.005 0 340.805 0.58 ;
 RECT 341.205 0 341.405 0.58 ;
 RECT 341.805 0 357.605 0.58 ;
 RECT 358.005 0 358.205 0.58 ;
 RECT 358.605 0 374.405 0.58 ;
 RECT 374.805 0 375.005 0.58 ;
 RECT 375.405 0 391.205 0.58 ;
 RECT 391.605 0 391.805 0.58 ;
 RECT 392.205 0 408.005 0.58 ;
 RECT 408.405 0 408.605 0.58 ;
 RECT 409.005 0 424.805 0.58 ;
 RECT 425.205 0 425.405 0.58 ;
 RECT 425.805 0 441.605 0.58 ;
 RECT 442.005 0 442.205 0.58 ;
 RECT 442.605 0 458.405 0.58 ;
 RECT 458.805 0 459.005 0.58 ;
 RECT 459.405 0 475.205 0.58 ;
 RECT 475.605 0 475.805 0.58 ;
 RECT 476.205 0 492.005 0.58 ;
 RECT 492.405 0 492.605 0.58 ;
 RECT 493.005 0 508.805 0.58 ;
 RECT 509.205 0 509.405 0.58 ;
 RECT 509.805 0 525.605 0.58 ;
 RECT 526.005 0 526.205 0.58 ;
 RECT 526.605 0 542.405 0.58 ;
 RECT 542.805 0 543.005 0.58 ;
 RECT 543.405 0 559.205 0.58 ;
 RECT 559.605 0 559.805 0.58 ;
 RECT 560.205 0 569.26 0.58 ;
 RECT 0 0.58 569.26 307.045 ;

 LAYER V1 ;
 RECT 0 0 569.26 307.045 ;
 LAYER V2 ;
 RECT 0 0 569.26 307.045 ;
 LAYER V3 ;
 RECT 0 0 569.26 307.045 ;

 LAYER M4 ;
 RECT 8.705 0 9.005 307.045 ;
 RECT 9.005 0 9.505 307.045 ;
 RECT 9.505 0 9.605 307.045 ;
 RECT 9.605 0 10.105 307.045 ;
 RECT 10.105 0 10.405 0.58 ;
 RECT 10.105 0.58 10.405 307.045 ;
 RECT 25.505 0 25.805 307.045 ;
 RECT 25.805 0 26.305 307.045 ;
 RECT 26.405 0 26.905 307.045 ;
 RECT 26.905 0 27.205 0.58 ;
 RECT 26.905 0.58 27.205 307.045 ;
 RECT 42.305 0 42.605 307.045 ;
 RECT 42.605 0 43.105 307.045 ;
 RECT 43.205 0 43.705 307.045 ;
 RECT 43.705 0 44.005 0.58 ;
 RECT 43.705 0.58 44.005 307.045 ;
 RECT 59.105 0 59.405 307.045 ;
 RECT 59.405 0 59.905 307.045 ;
 RECT 59.905 0 60.005 307.045 ;
 RECT 60.005 0 60.505 307.045 ;
 RECT 60.505 0 60.805 0.58 ;
 RECT 60.505 0.58 60.805 307.045 ;
 RECT 75.905 0 76.205 307.045 ;
 RECT 76.205 0 76.705 307.045 ;
 RECT 76.705 0 76.805 307.045 ;
 RECT 76.805 0 77.305 307.045 ;
 RECT 77.305 0 77.605 0.58 ;
 RECT 77.305 0.58 77.605 307.045 ;
 RECT 92.705 0 93.005 307.045 ;
 RECT 93.005 0 93.505 307.045 ;
 RECT 93.605 0 94.105 307.045 ;
 RECT 94.105 0 94.405 0.58 ;
 RECT 94.105 0.58 94.405 307.045 ;
 RECT 109.505 0 109.805 307.045 ;
 RECT 109.805 0 110.305 307.045 ;
 RECT 110.405 0 110.905 307.045 ;
 RECT 110.905 0 111.205 0.58 ;
 RECT 110.905 0.58 111.205 307.045 ;
 RECT 126.305 0 126.605 307.045 ;
 RECT 126.605 0 127.105 307.045 ;
 RECT 127.205 0 127.705 307.045 ;
 RECT 127.705 0 128.005 0.58 ;
 RECT 127.705 0.58 128.005 307.045 ;
 RECT 143.105 0 143.405 307.045 ;
 RECT 143.405 0 143.905 307.045 ;
 RECT 143.905 0 144.005 307.045 ;
 RECT 144.005 0 144.505 307.045 ;
 RECT 144.505 0 144.805 0.58 ;
 RECT 144.505 0.58 144.805 307.045 ;
 RECT 159.905 0 160.205 307.045 ;
 RECT 160.205 0 160.705 307.045 ;
 RECT 160.705 0 160.805 307.045 ;
 RECT 160.805 0 161.305 307.045 ;
 RECT 161.305 0 161.605 0.58 ;
 RECT 161.305 0.58 161.605 307.045 ;
 RECT 176.705 0 177.005 307.045 ;
 RECT 177.005 0 177.505 307.045 ;
 RECT 177.605 0 178.105 307.045 ;
 RECT 178.105 0 178.405 0.58 ;
 RECT 178.105 0.58 178.405 307.045 ;
 RECT 193.505 0 193.805 307.045 ;
 RECT 193.805 0 194.305 307.045 ;
 RECT 194.405 0 194.905 307.045 ;
 RECT 194.905 0 195.205 0.58 ;
 RECT 194.905 0.58 195.205 307.045 ;
 RECT 210.305 0 210.605 307.045 ;
 RECT 210.605 0 211.105 307.045 ;
 RECT 211.205 0 211.705 307.045 ;
 RECT 211.705 0 212.005 0.58 ;
 RECT 211.705 0.58 212.005 307.045 ;
 RECT 227.105 0 227.405 307.045 ;
 RECT 227.405 0 227.905 307.045 ;
 RECT 227.905 0 228.005 307.045 ;
 RECT 228.005 0 228.505 307.045 ;
 RECT 228.505 0 228.805 0.58 ;
 RECT 228.505 0.58 228.805 307.045 ;
 RECT 243.905 0 244.205 307.045 ;
 RECT 244.205 0 244.705 307.045 ;
 RECT 244.705 0 244.805 307.045 ;
 RECT 244.805 0 245.305 307.045 ;
 RECT 245.305 0 245.605 0.58 ;
 RECT 245.305 0.58 245.605 307.045 ;
 RECT 260.705 0 261.005 307.045 ;
 RECT 261.005 0 261.505 307.045 ;
 RECT 261.605 0 262.105 307.045 ;
 RECT 262.105 0 262.405 0.58 ;
 RECT 262.105 0.58 262.405 307.045 ;
 RECT 269.105 0 270.325 307.045 ;
 RECT 270.325 0 270.725 307.045 ;
 RECT 270.725 0 271.125 307.045 ;
 RECT 271.125 0 271.525 307.045 ;
 RECT 271.525 0 272.205 0.58 ;
 RECT 271.525 0.58 272.205 307.045 ;
 RECT 274.305 0 274.505 0.58 ;
 RECT 274.305 0.58 274.505 307.045 ;
 RECT 274.305 0 274.505 307.045 ;
 RECT 276.605 0 277.205 307.045 ;
 RECT 277.205 0 277.605 307.045 ;
 RECT 277.605 0 277.805 0.58 ;
 RECT 277.605 0.58 277.805 307.045 ;
 RECT 279.905 0 280.505 307.045 ;
 RECT 280.505 0 280.955 307.045 ;
 RECT 280.955 0 281.405 307.045 ;
 RECT 281.405 0 281.855 307.045 ;
 RECT 281.855 0 282.31 307.045 ;
 RECT 282.31 0 283.495 0.58 ;
 RECT 282.31 0.58 283.495 307.045 ;
 RECT 285.695 0 285.895 0.58 ;
 RECT 285.695 0.58 285.895 307.045 ;
 RECT 285.695 0 285.895 307.045 ;
 RECT 288.095 0 288.695 307.045 ;
 RECT 288.695 0 289.095 307.045 ;
 RECT 289.095 0 289.495 307.045 ;
 RECT 289.495 0 289.695 0.58 ;
 RECT 289.495 0.58 289.695 307.045 ;
 RECT 291.895 0 292.48 307.045 ;
 RECT 292.48 0 292.68 0.58 ;
 RECT 292.48 0.58 292.68 307.045 ;
 RECT 294.88 0 295.08 0.58 ;
 RECT 294.88 0.58 295.08 307.045 ;
 RECT 294.88 0 295.08 307.045 ;
 RECT 297.28 0 298.495 307.045 ;
 RECT 298.495 0 300.155 0.58 ;
 RECT 298.495 0.58 300.155 307.045 ;
 RECT 306.855 0 307.155 307.045 ;
 RECT 307.155 0 307.655 307.045 ;
 RECT 307.755 0 308.255 307.045 ;
 RECT 308.255 0 308.555 0.58 ;
 RECT 308.255 0.58 308.555 307.045 ;
 RECT 323.655 0 323.955 307.045 ;
 RECT 323.955 0 324.455 307.045 ;
 RECT 324.455 0 324.555 307.045 ;
 RECT 324.555 0 325.055 307.045 ;
 RECT 325.055 0 325.355 0.58 ;
 RECT 325.055 0.58 325.355 307.045 ;
 RECT 340.455 0 340.755 307.045 ;
 RECT 340.755 0 341.255 307.045 ;
 RECT 341.255 0 341.355 307.045 ;
 RECT 341.355 0 341.855 307.045 ;
 RECT 341.855 0 342.155 0.58 ;
 RECT 341.855 0.58 342.155 307.045 ;
 RECT 357.255 0 357.555 307.045 ;
 RECT 357.555 0 358.055 307.045 ;
 RECT 358.055 0 358.155 307.045 ;
 RECT 358.155 0 358.655 307.045 ;
 RECT 358.655 0 358.955 0.58 ;
 RECT 358.655 0.58 358.955 307.045 ;
 RECT 374.055 0 374.355 307.045 ;
 RECT 374.355 0 374.855 307.045 ;
 RECT 374.855 0 374.955 307.045 ;
 RECT 374.955 0 375.455 307.045 ;
 RECT 375.455 0 375.755 0.58 ;
 RECT 375.455 0.58 375.755 307.045 ;
 RECT 390.855 0 391.155 307.045 ;
 RECT 391.155 0 391.655 307.045 ;
 RECT 391.755 0 392.255 307.045 ;
 RECT 392.255 0 392.555 0.58 ;
 RECT 392.255 0.58 392.555 307.045 ;
 RECT 407.655 0 407.955 307.045 ;
 RECT 407.955 0 408.455 307.045 ;
 RECT 408.555 0 409.055 307.045 ;
 RECT 409.055 0 409.355 0.58 ;
 RECT 409.055 0.58 409.355 307.045 ;
 RECT 424.455 0 424.755 307.045 ;
 RECT 424.755 0 425.255 307.045 ;
 RECT 425.255 0 425.355 307.045 ;
 RECT 425.355 0 425.855 307.045 ;
 RECT 425.855 0 426.155 0.58 ;
 RECT 425.855 0.58 426.155 307.045 ;
 RECT 441.255 0 441.555 307.045 ;
 RECT 441.555 0 442.055 307.045 ;
 RECT 442.055 0 442.155 307.045 ;
 RECT 442.155 0 442.655 307.045 ;
 RECT 442.655 0 442.955 0.58 ;
 RECT 442.655 0.58 442.955 307.045 ;
 RECT 458.055 0 458.355 307.045 ;
 RECT 458.355 0 458.855 307.045 ;
 RECT 458.855 0 458.955 307.045 ;
 RECT 458.955 0 459.455 307.045 ;
 RECT 459.455 0 459.755 0.58 ;
 RECT 459.455 0.58 459.755 307.045 ;
 RECT 474.855 0 475.155 307.045 ;
 RECT 475.155 0 475.655 307.045 ;
 RECT 475.655 0 475.755 307.045 ;
 RECT 475.755 0 476.255 307.045 ;
 RECT 476.255 0 476.555 0.58 ;
 RECT 476.255 0.58 476.555 307.045 ;
 RECT 491.655 0 491.955 307.045 ;
 RECT 491.955 0 492.455 307.045 ;
 RECT 492.555 0 493.055 307.045 ;
 RECT 493.055 0 493.355 0.58 ;
 RECT 493.055 0.58 493.355 307.045 ;
 RECT 508.455 0 508.755 307.045 ;
 RECT 508.755 0 509.255 307.045 ;
 RECT 509.255 0 509.355 307.045 ;
 RECT 509.355 0 509.855 307.045 ;
 RECT 509.855 0 510.155 0.58 ;
 RECT 509.855 0.58 510.155 307.045 ;
 RECT 525.255 0 525.555 307.045 ;
 RECT 525.555 0 526.055 307.045 ;
 RECT 526.155 0 526.655 307.045 ;
 RECT 526.655 0 526.955 0.58 ;
 RECT 526.655 0.58 526.955 307.045 ;
 RECT 542.055 0 542.355 307.045 ;
 RECT 542.355 0 542.855 307.045 ;
 RECT 542.855 0 542.955 307.045 ;
 RECT 542.955 0 543.455 307.045 ;
 RECT 543.455 0 543.755 0.58 ;
 RECT 543.455 0.58 543.755 307.045 ;
 RECT 558.855 0 559.155 307.045 ;
 RECT 559.155 0 559.655 307.045 ;
 RECT 559.655 0 559.755 307.045 ;
 RECT 559.755 0 560.255 307.045 ;
 RECT 560.255 0 560.555 0.58 ;
 RECT 560.255 0.58 560.555 307.045 ;
 LAYER V4 ;
 RECT 8.705 0 9.005 307.045 ;
 RECT 9.005 0 9.505 307.045 ;
 RECT 9.505 0 9.605 307.045 ;
 RECT 9.605 0 10.105 307.045 ;
 RECT 10.105 0 10.405 0.58 ;
 RECT 10.105 0.58 10.405 307.045 ;
 RECT 25.505 0 25.805 307.045 ;
 RECT 25.805 0 26.305 307.045 ;
 RECT 26.405 0 26.905 307.045 ;
 RECT 26.905 0 27.205 0.58 ;
 RECT 26.905 0.58 27.205 307.045 ;
 RECT 42.305 0 42.605 307.045 ;
 RECT 42.605 0 43.105 307.045 ;
 RECT 43.205 0 43.705 307.045 ;
 RECT 43.705 0 44.005 0.58 ;
 RECT 43.705 0.58 44.005 307.045 ;
 RECT 59.105 0 59.405 307.045 ;
 RECT 59.405 0 59.905 307.045 ;
 RECT 59.905 0 60.005 307.045 ;
 RECT 60.005 0 60.505 307.045 ;
 RECT 60.505 0 60.805 0.58 ;
 RECT 60.505 0.58 60.805 307.045 ;
 RECT 75.905 0 76.205 307.045 ;
 RECT 76.205 0 76.705 307.045 ;
 RECT 76.705 0 76.805 307.045 ;
 RECT 76.805 0 77.305 307.045 ;
 RECT 77.305 0 77.605 0.58 ;
 RECT 77.305 0.58 77.605 307.045 ;
 RECT 92.705 0 93.005 307.045 ;
 RECT 93.005 0 93.505 307.045 ;
 RECT 93.605 0 94.105 307.045 ;
 RECT 94.105 0 94.405 0.58 ;
 RECT 94.105 0.58 94.405 307.045 ;
 RECT 109.505 0 109.805 307.045 ;
 RECT 109.805 0 110.305 307.045 ;
 RECT 110.405 0 110.905 307.045 ;
 RECT 110.905 0 111.205 0.58 ;
 RECT 110.905 0.58 111.205 307.045 ;
 RECT 126.305 0 126.605 307.045 ;
 RECT 126.605 0 127.105 307.045 ;
 RECT 127.205 0 127.705 307.045 ;
 RECT 127.705 0 128.005 0.58 ;
 RECT 127.705 0.58 128.005 307.045 ;
 RECT 143.105 0 143.405 307.045 ;
 RECT 143.405 0 143.905 307.045 ;
 RECT 143.905 0 144.005 307.045 ;
 RECT 144.005 0 144.505 307.045 ;
 RECT 144.505 0 144.805 0.58 ;
 RECT 144.505 0.58 144.805 307.045 ;
 RECT 159.905 0 160.205 307.045 ;
 RECT 160.205 0 160.705 307.045 ;
 RECT 160.705 0 160.805 307.045 ;
 RECT 160.805 0 161.305 307.045 ;
 RECT 161.305 0 161.605 0.58 ;
 RECT 161.305 0.58 161.605 307.045 ;
 RECT 176.705 0 177.005 307.045 ;
 RECT 177.005 0 177.505 307.045 ;
 RECT 177.605 0 178.105 307.045 ;
 RECT 178.105 0 178.405 0.58 ;
 RECT 178.105 0.58 178.405 307.045 ;
 RECT 193.505 0 193.805 307.045 ;
 RECT 193.805 0 194.305 307.045 ;
 RECT 194.405 0 194.905 307.045 ;
 RECT 194.905 0 195.205 0.58 ;
 RECT 194.905 0.58 195.205 307.045 ;
 RECT 210.305 0 210.605 307.045 ;
 RECT 210.605 0 211.105 307.045 ;
 RECT 211.205 0 211.705 307.045 ;
 RECT 211.705 0 212.005 0.58 ;
 RECT 211.705 0.58 212.005 307.045 ;
 RECT 227.105 0 227.405 307.045 ;
 RECT 227.405 0 227.905 307.045 ;
 RECT 227.905 0 228.005 307.045 ;
 RECT 228.005 0 228.505 307.045 ;
 RECT 228.505 0 228.805 0.58 ;
 RECT 228.505 0.58 228.805 307.045 ;
 RECT 243.905 0 244.205 307.045 ;
 RECT 244.205 0 244.705 307.045 ;
 RECT 244.705 0 244.805 307.045 ;
 RECT 244.805 0 245.305 307.045 ;
 RECT 245.305 0 245.605 0.58 ;
 RECT 245.305 0.58 245.605 307.045 ;
 RECT 260.705 0 261.005 307.045 ;
 RECT 261.005 0 261.505 307.045 ;
 RECT 261.605 0 262.105 307.045 ;
 RECT 262.105 0 262.405 0.58 ;
 RECT 262.105 0.58 262.405 307.045 ;
 RECT 269.105 0 270.325 307.045 ;
 RECT 270.325 0 270.725 307.045 ;
 RECT 270.725 0 271.125 307.045 ;
 RECT 271.125 0 271.525 307.045 ;
 RECT 271.525 0 272.205 0.58 ;
 RECT 271.525 0.58 272.205 307.045 ;
 RECT 274.305 0 274.505 0.58 ;
 RECT 274.305 0.58 274.505 307.045 ;
 RECT 274.305 0 274.505 307.045 ;
 RECT 276.605 0 277.205 307.045 ;
 RECT 277.205 0 277.605 307.045 ;
 RECT 277.605 0 277.805 0.58 ;
 RECT 277.605 0.58 277.805 307.045 ;
 RECT 279.905 0 280.505 307.045 ;
 RECT 280.505 0 280.955 307.045 ;
 RECT 280.955 0 281.405 307.045 ;
 RECT 281.405 0 281.855 307.045 ;
 RECT 281.855 0 282.31 307.045 ;
 RECT 282.31 0 283.495 0.58 ;
 RECT 282.31 0.58 283.495 307.045 ;
 RECT 285.695 0 285.895 0.58 ;
 RECT 285.695 0.58 285.895 307.045 ;
 RECT 285.695 0 285.895 307.045 ;
 RECT 288.095 0 288.695 307.045 ;
 RECT 288.695 0 289.095 307.045 ;
 RECT 289.095 0 289.495 307.045 ;
 RECT 289.495 0 289.695 0.58 ;
 RECT 289.495 0.58 289.695 307.045 ;
 RECT 291.895 0 292.48 307.045 ;
 RECT 292.48 0 292.68 0.58 ;
 RECT 292.48 0.58 292.68 307.045 ;
 RECT 294.88 0 295.08 0.58 ;
 RECT 294.88 0.58 295.08 307.045 ;
 RECT 294.88 0 295.08 307.045 ;
 RECT 297.28 0 298.495 307.045 ;
 RECT 298.495 0 300.155 0.58 ;
 RECT 298.495 0.58 300.155 307.045 ;
 RECT 306.855 0 307.155 307.045 ;
 RECT 307.155 0 307.655 307.045 ;
 RECT 307.755 0 308.255 307.045 ;
 RECT 308.255 0 308.555 0.58 ;
 RECT 308.255 0.58 308.555 307.045 ;
 RECT 323.655 0 323.955 307.045 ;
 RECT 323.955 0 324.455 307.045 ;
 RECT 324.455 0 324.555 307.045 ;
 RECT 324.555 0 325.055 307.045 ;
 RECT 325.055 0 325.355 0.58 ;
 RECT 325.055 0.58 325.355 307.045 ;
 RECT 340.455 0 340.755 307.045 ;
 RECT 340.755 0 341.255 307.045 ;
 RECT 341.255 0 341.355 307.045 ;
 RECT 341.355 0 341.855 307.045 ;
 RECT 341.855 0 342.155 0.58 ;
 RECT 341.855 0.58 342.155 307.045 ;
 RECT 357.255 0 357.555 307.045 ;
 RECT 357.555 0 358.055 307.045 ;
 RECT 358.055 0 358.155 307.045 ;
 RECT 358.155 0 358.655 307.045 ;
 RECT 358.655 0 358.955 0.58 ;
 RECT 358.655 0.58 358.955 307.045 ;
 RECT 374.055 0 374.355 307.045 ;
 RECT 374.355 0 374.855 307.045 ;
 RECT 374.855 0 374.955 307.045 ;
 RECT 374.955 0 375.455 307.045 ;
 RECT 375.455 0 375.755 0.58 ;
 RECT 375.455 0.58 375.755 307.045 ;
 RECT 390.855 0 391.155 307.045 ;
 RECT 391.155 0 391.655 307.045 ;
 RECT 391.755 0 392.255 307.045 ;
 RECT 392.255 0 392.555 0.58 ;
 RECT 392.255 0.58 392.555 307.045 ;
 RECT 407.655 0 407.955 307.045 ;
 RECT 407.955 0 408.455 307.045 ;
 RECT 408.555 0 409.055 307.045 ;
 RECT 409.055 0 409.355 0.58 ;
 RECT 409.055 0.58 409.355 307.045 ;
 RECT 424.455 0 424.755 307.045 ;
 RECT 424.755 0 425.255 307.045 ;
 RECT 425.255 0 425.355 307.045 ;
 RECT 425.355 0 425.855 307.045 ;
 RECT 425.855 0 426.155 0.58 ;
 RECT 425.855 0.58 426.155 307.045 ;
 RECT 441.255 0 441.555 307.045 ;
 RECT 441.555 0 442.055 307.045 ;
 RECT 442.055 0 442.155 307.045 ;
 RECT 442.155 0 442.655 307.045 ;
 RECT 442.655 0 442.955 0.58 ;
 RECT 442.655 0.58 442.955 307.045 ;
 RECT 458.055 0 458.355 307.045 ;
 RECT 458.355 0 458.855 307.045 ;
 RECT 458.855 0 458.955 307.045 ;
 RECT 458.955 0 459.455 307.045 ;
 RECT 459.455 0 459.755 0.58 ;
 RECT 459.455 0.58 459.755 307.045 ;
 RECT 474.855 0 475.155 307.045 ;
 RECT 475.155 0 475.655 307.045 ;
 RECT 475.655 0 475.755 307.045 ;
 RECT 475.755 0 476.255 307.045 ;
 RECT 476.255 0 476.555 0.58 ;
 RECT 476.255 0.58 476.555 307.045 ;
 RECT 491.655 0 491.955 307.045 ;
 RECT 491.955 0 492.455 307.045 ;
 RECT 492.555 0 493.055 307.045 ;
 RECT 493.055 0 493.355 0.58 ;
 RECT 493.055 0.58 493.355 307.045 ;
 RECT 508.455 0 508.755 307.045 ;
 RECT 508.755 0 509.255 307.045 ;
 RECT 509.255 0 509.355 307.045 ;
 RECT 509.355 0 509.855 307.045 ;
 RECT 509.855 0 510.155 0.58 ;
 RECT 509.855 0.58 510.155 307.045 ;
 RECT 525.255 0 525.555 307.045 ;
 RECT 525.555 0 526.055 307.045 ;
 RECT 526.155 0 526.655 307.045 ;
 RECT 526.655 0 526.955 0.58 ;
 RECT 526.655 0.58 526.955 307.045 ;
 RECT 542.055 0 542.355 307.045 ;
 RECT 542.355 0 542.855 307.045 ;
 RECT 542.855 0 542.955 307.045 ;
 RECT 542.955 0 543.455 307.045 ;
 RECT 543.455 0 543.755 0.58 ;
 RECT 543.455 0.58 543.755 307.045 ;
 RECT 558.855 0 559.155 307.045 ;
 RECT 559.155 0 559.655 307.045 ;
 RECT 559.655 0 559.755 307.045 ;
 RECT 559.755 0 560.255 307.045 ;
 RECT 560.255 0 560.555 0.58 ;
 RECT 560.255 0.58 560.555 307.045 ;
 END

END S55NLLGSPH_X512Y16D32
END LIBRARY