************************************************************************
* auCdl Netlist:
*
* Library Name:  SMIC_MEMORY
* Top Cell Name: S55NLLGSPH_X512Y16D32
* Version:  V1.1
* View Name:     schematic
* Netlisted on:  Wed Feb 15 21:09:21 CST 2023
************************************************************************
*.BIPOLAR
*.RESI = 2000
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM


************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_BLSTRAP1
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_BLSTRAP1 BL VDD VSS
MN1 BL VSS NET21 VSS STNPGHVT W=85.000N L=75.00N M=1
MN0 NET18 VSS VSS VSS STNPDHVT W=135.000N L=65.000N M=1
MP0 NET26 VSS VDD VDD STPLHVT W=85.000N L=65.000N M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP B BX VDD VSS WL1
MTA1 BX VSS NET37 VSS STNPGHVT W=85.000N L=75.00N M=1
MTA0 B WL1 NET46 VSS STNPGHVT W=85.000N L=75.00N M=1
MTD1 NET37 NET46 VSS VSS STNPDHVT W=135.000N L=65.000N M=1
MTD0 NET46 NET37 VSS VSS STNPDHVT W=135.000N L=65.000N M=1
MTL1 NET37 NET46 VDD VDD STPLHVT W=85.000N L=65.000N M=1
MTL0 NET46 NET37 VDD VDD STPLHVT W=85.000N L=65.000N M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP4B
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP4B BX0 BX1 VDD VSS WL[3] WL[2] WL[1] WL[0]
XI5 NET29 BX1 VDD VSS WL[3] S55NLLGSPH_X512Y16D32_PCAP
XI4 NET29 NET32 VDD VSS WL[2] S55NLLGSPH_X512Y16D32_PCAP
XI3 NET39 NET32 VDD VSS WL[1] S55NLLGSPH_X512Y16D32_PCAP
XI2 NET39 BX0 VDD VSS WL[0] S55NLLGSPH_X512Y16D32_PCAP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP64B
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP64B B0 B1 VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XI0 NET31 NET61 VDD VSS WL[7] WL[6] WL[5] WL[4] S55NLLGSPH_X512Y16D32_PCAP4B
XI1 B0 NET31 VDD VSS WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_PCAP4B
XI2 NET01 NET32 VDD VSS WL[11] WL[10] WL[9] WL[8] S55NLLGSPH_X512Y16D32_PCAP4B
XI3 NET32 NET61 VDD VSS WL[15] WL[14] WL[13] WL[12] S55NLLGSPH_X512Y16D32_PCAP4B
XI4 NET33 NET62 VDD VSS WL[23] WL[22] WL[21] WL[20] S55NLLGSPH_X512Y16D32_PCAP4B
XI5 NET01 NET33 VDD VSS WL[19] WL[18] WL[17] WL[16] S55NLLGSPH_X512Y16D32_PCAP4B
XI6 NET02 NET34 VDD VSS WL[27] WL[26] WL[25] WL[24] S55NLLGSPH_X512Y16D32_PCAP4B
XI7 NET34 NET62 VDD VSS WL[31] WL[30] WL[29] WL[28] S55NLLGSPH_X512Y16D32_PCAP4B
XI8 NET35 NET63 VDD VSS WL[39] WL[38] WL[37] WL[36] S55NLLGSPH_X512Y16D32_PCAP4B
XI9 NET02 NET35 VDD VSS WL[35] WL[34] WL[33] WL[32] S55NLLGSPH_X512Y16D32_PCAP4B
XI10 NET03 NET36 VDD VSS WL[43] WL[42] WL[41] WL[40] S55NLLGSPH_X512Y16D32_PCAP4B
XI11 NET36 NET63 VDD VSS WL[47] WL[46] WL[45] WL[44] S55NLLGSPH_X512Y16D32_PCAP4B
XI12 NET37 NET64 VDD VSS WL[55] WL[54] WL[53] WL[52] S55NLLGSPH_X512Y16D32_PCAP4B
XI13 NET03 NET37 VDD VSS WL[51] WL[50] WL[49] WL[48] S55NLLGSPH_X512Y16D32_PCAP4B
XI14 B1 NET38 VDD VSS WL[59] WL[58] WL[57] WL[56] S55NLLGSPH_X512Y16D32_PCAP4B
XI15 NET38 NET64 VDD VSS WL[63] WL[62] WL[61] WL[60] S55NLLGSPH_X512Y16D32_PCAP4B
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP_EDGE66B_RED
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP_EDGE66B_RED RWL0 RWL1 VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XI0 NET44 VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI1 NET48 NET44 VDD VSS RWL0 S55NLLGSPH_X512Y16D32_PCAP
XI2 NET48 NET49 VDD VSS RWL1 S55NLLGSPH_X512Y16D32_PCAP
XI3 NET49 NET36 VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_PCAP64B
XI4 NET36 VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP4A
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP4A B0 B1 VDD VSS WL[3] WL[2] WL[1] WL[0]
XI5 B1 NET27 VDD VSS WL[3] S55NLLGSPH_X512Y16D32_PCAP
XI4 NET34 NET27 VDD VSS WL[2] S55NLLGSPH_X512Y16D32_PCAP
XI3 NET34 NET37 VDD VSS WL[1] S55NLLGSPH_X512Y16D32_PCAP
XI2 B0 NET37 VDD VSS WL[0] S55NLLGSPH_X512Y16D32_PCAP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP64A
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP64A B0 B1 VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XI0 NET31 NET61 VDD VSS WL[7] WL[6] WL[5] WL[4] S55NLLGSPH_X512Y16D32_PCAP4A
XI1 B0 NET31 VDD VSS WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_PCAP4A
XI2 NET01 NET32 VDD VSS WL[11] WL[10] WL[9] WL[8] S55NLLGSPH_X512Y16D32_PCAP4A
XI3 NET32 NET61 VDD VSS WL[15] WL[14] WL[13] WL[12] S55NLLGSPH_X512Y16D32_PCAP4A
XI4 NET33 NET62 VDD VSS WL[23] WL[22] WL[21] WL[20] S55NLLGSPH_X512Y16D32_PCAP4A
XI5 NET01 NET33 VDD VSS WL[19] WL[18] WL[17] WL[16] S55NLLGSPH_X512Y16D32_PCAP4A
XI6 NET02 NET34 VDD VSS WL[27] WL[26] WL[25] WL[24] S55NLLGSPH_X512Y16D32_PCAP4A
XI7 NET34 NET62 VDD VSS WL[31] WL[30] WL[29] WL[28] S55NLLGSPH_X512Y16D32_PCAP4A
XI8 NET35 NET63 VDD VSS WL[39] WL[38] WL[37] WL[36] S55NLLGSPH_X512Y16D32_PCAP4A
XI9 NET02 NET35 VDD VSS WL[35] WL[34] WL[33] WL[32] S55NLLGSPH_X512Y16D32_PCAP4A
XI10 NET03 NET36 VDD VSS WL[43] WL[42] WL[41] WL[40] S55NLLGSPH_X512Y16D32_PCAP4A
XI11 NET36 NET63 VDD VSS WL[47] WL[46] WL[45] WL[44] S55NLLGSPH_X512Y16D32_PCAP4A
XI12 NET37 NET64 VDD VSS WL[55] WL[54] WL[53] WL[52] S55NLLGSPH_X512Y16D32_PCAP4A
XI13 NET03 NET37 VDD VSS WL[51] WL[50] WL[49] WL[48] S55NLLGSPH_X512Y16D32_PCAP4A
XI14 B1 NET38 VDD VSS WL[59] WL[58] WL[57] WL[56] S55NLLGSPH_X512Y16D32_PCAP4A
XI15 NET38 NET64 VDD VSS WL[63] WL[62] WL[61] WL[60] S55NLLGSPH_X512Y16D32_PCAP4A
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP_EDGE64A
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP_EDGE64A VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XI0 NET49 VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI1 NET49 NET36 VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_PCAP64A
XI2 NET36 VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP_EDGE64B
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP_EDGE64B VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XI0 NET49 VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI1 NET49 NET36 VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_PCAP64B
XI2 NET36 VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP4B_RDWL
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP4B_RDWL BX0 BX1 VDD VSS WL[0] WL[1] WL[2] WL[3]
XI5 NET29 BX1 VDD VSS WL[3] S55NLLGSPH_X512Y16D32_PCAP
XI4 NET29 NET32 VDD VSS WL[2] S55NLLGSPH_X512Y16D32_PCAP
XI3 NET39 NET32 VDD VSS WL[1] S55NLLGSPH_X512Y16D32_PCAP
XI2 NET39 BX0 VDD VSS WL[0] S55NLLGSPH_X512Y16D32_PCAP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP_EDGE68A_TOP
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP_EDGE68A_TOP STWL VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57]
+WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47]
+WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37]
+WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27]
+WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17]
+WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7]
+WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XI0 NET49 VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI1 NET49 NET36 VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_PCAP64A
XI2 NET36 NET40 VDD VSS VSS STWL STWL VSS S55NLLGSPH_X512Y16D32_PCAP4B_RDWL
XI3 NET40 VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP_EDGE256_DOWN
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP_EDGE256_DOWN RWL0 RWL1 STWL VDD VSS WL[255] WL[254] WL[253] WL[252] WL[251]
+WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241]
+WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231]
+WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221]
+WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211]
+WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201]
+WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191]
+WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181]
+WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171]
+WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161]
+WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151]
+WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141]
+WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131]
+WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121]
+WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111]
+WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101]
+WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91]
+WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81]
+WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71]
+WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61]
+WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51]
+WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41]
+WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31]
+WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21]
+WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11]
+WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1]
+WL[0]
XI0 RWL0 RWL1 VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_PCAP_EDGE66B_RED
XI1 VDD VSS WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120]
+WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110]
+WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100]
+WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90]
+WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80]
+WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70]
+WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] S55NLLGSPH_X512Y16D32_PCAP_EDGE64A
XI2 VDD VSS WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184]
+WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174]
+WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164]
+WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154]
+WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144]
+WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134]
+WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] S55NLLGSPH_X512Y16D32_PCAP_EDGE64B
XI3 STWL VDD VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249]
+WL[248] WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239]
+WL[238] WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229]
+WL[228] WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219]
+WL[218] WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209]
+WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199]
+WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] S55NLLGSPH_X512Y16D32_PCAP_EDGE68A_TOP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525 B BX VDD VSS WL1
MM2 BX WL1 BCN VSS STNPGHVT W=85.000N L=75.00N M=1
MM3 B WL1 BC VSS STNPGHVT W=85.000N L=75.00N M=1
MM0 BCN BC VSS VSS STNPDHVT W=135.00N L=65.00N M=1
MM1 BC BCN VSS VSS STNPDHVT W=135.00N L=65.00N M=1
MM5 BCN BC VDD VDD STPLHVT W=85.000N L=65.00N M=1
MM6 BC BCN VDD VDD STPLHVT W=85.000N L=65.00N M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_BITCELL2X2
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_BITCELL2X2 B[1] B[0] BX[1] BX[0] VDD VSS WL[1] WL[0]
XI8 B[1] BX[1] VDD VSS WL[1] S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525
XI9 B[0] BX[0] VDD VSS WL[1] S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525
XI7 B[1] BX[1] VDD VSS WL[0] S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525
XI5 B[0] BX[0] VDD VSS WL[0] S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_BITCELLREDUNDANCE2X2
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_BITCELLREDUNDANCE2X2 B[1] B[0] BX[1] BX[0] RWL[0] RWL[1] VDD VSS
XI8 B[1] BX[1] VDD VSS RWL[1] S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525
XI9 B[0] BX[0] VDD VSS RWL[1] S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525
XI7 B[1] BX[1] VDD VSS RWL[0] S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525
XI5 B[0] BX[0] VDD VSS RWL[0] S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_BITCELL66X2A_RED
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_BITCELL66X2A_RED BL[1] BL[0] BLX[1] BLX[0] RWL[0] RWL[1] VDD VSS WL[63] WL[62]
+WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52]
+WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42]
+WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32]
+WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22]
+WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12]
+WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2]
+WL[1] WL[0]
XI0 BLX[1] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI1 BLX[0] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI2 BLX[1] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI3 BLX[0] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI4 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI5 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[3] WL[2] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI6 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[5] WL[4] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI7 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[7] WL[6] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI8 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[9] WL[8] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI9 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[11] WL[10] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI10 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[13] WL[12] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI11 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[15] WL[14] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI12 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[17] WL[16] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI13 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[19] WL[18] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI14 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[21] WL[20] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI15 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[23] WL[22] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI16 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[25] WL[24] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI17 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[27] WL[26] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI18 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[29] WL[28] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI19 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[31] WL[30] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI20 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[33] WL[32] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI21 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[35] WL[34] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI22 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[37] WL[36] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI23 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[39] WL[38] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI24 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[41] WL[40] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI25 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[43] WL[42] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI26 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[45] WL[44] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI27 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[47] WL[46] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI28 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[49] WL[48] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI29 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[51] WL[50] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI30 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[53] WL[52] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI31 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[55] WL[54] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI32 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[57] WL[56] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI33 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[59] WL[58] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI34 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[61] WL[60] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI35 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[63] WL[62] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI36 BL[1] BL[0] BLX[1] BLX[0] RWL[0] RWL[1] VDD VSS S55NLLGSPH_X512Y16D32_BITCELLREDUNDANCE2X2
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_BITCELL64X2B
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_BITCELL64X2B BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[63] WL[62] WL[61] WL[60]
+WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50]
+WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40]
+WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30]
+WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20]
+WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10]
+WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XI0 BL[1] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI1 BL[0] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI2 BL[1] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI3 BL[0] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI4 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI5 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[3] WL[2] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI6 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[5] WL[4] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI7 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[7] WL[6] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI8 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[9] WL[8] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI9 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[11] WL[10] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI10 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[13] WL[12] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI11 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[15] WL[14] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI12 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[17] WL[16] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI13 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[19] WL[18] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI14 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[21] WL[20] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI15 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[23] WL[22] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI16 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[25] WL[24] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI17 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[27] WL[26] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI18 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[29] WL[28] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI19 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[31] WL[30] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI20 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[33] WL[32] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI21 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[35] WL[34] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI22 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[37] WL[36] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI23 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[39] WL[38] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI24 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[41] WL[40] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI25 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[43] WL[42] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI26 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[45] WL[44] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI27 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[47] WL[46] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI28 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[49] WL[48] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI29 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[51] WL[50] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI30 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[53] WL[52] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI31 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[55] WL[54] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI32 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[57] WL[56] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI33 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[59] WL[58] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI34 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[61] WL[60] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI35 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[63] WL[62] S55NLLGSPH_X512Y16D32_BITCELL2X2
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_BITCELL64X2A
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_BITCELL64X2A BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[63] WL[62] WL[61] WL[60]
+WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50]
+WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40]
+WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30]
+WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20]
+WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10]
+WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XI0 BLX[1] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI1 BLX[0] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI2 BLX[1] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI3 BLX[0] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI4 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI5 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[3] WL[2] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI6 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[5] WL[4] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI7 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[7] WL[6] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI8 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[9] WL[8] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI9 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[11] WL[10] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI10 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[13] WL[12] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI11 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[15] WL[14] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI12 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[17] WL[16] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI13 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[19] WL[18] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI14 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[21] WL[20] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI15 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[23] WL[22] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI16 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[25] WL[24] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI17 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[27] WL[26] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI18 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[29] WL[28] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI19 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[31] WL[30] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI20 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[33] WL[32] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI21 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[35] WL[34] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI22 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[37] WL[36] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI23 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[39] WL[38] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI24 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[41] WL[40] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI25 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[43] WL[42] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI26 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[45] WL[44] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI27 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[47] WL[46] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI28 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[49] WL[48] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI29 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[51] WL[50] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI30 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[53] WL[52] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI31 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[55] WL[54] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI32 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[57] WL[56] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI33 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[59] WL[58] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI34 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[61] WL[60] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI35 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[63] WL[62] S55NLLGSPH_X512Y16D32_BITCELL2X2
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_BITCELL_RDWL2B
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_BITCELL_RDWL2B BL0 BL1 VDD VSS WL0 WL1
XI5 BL0 NET11 VDD VSS WL0 S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525
XI6 BL1 NET11 VDD VSS WL1 S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_BITCELL68X2B_TOP
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_BITCELL68X2B_TOP BL[1] BL[0] BLX[1] BLX[0] RDWL VDD VSS WL[63] WL[62] WL[61]
+WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51]
+WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41]
+WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31]
+WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21]
+WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11]
+WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1]
+WL[0]
XI0 BL[0] NET44[1] VDD VSS VSS RDWL S55NLLGSPH_X512Y16D32_BITCELL_RDWL2B
XI1 BL[1] NET44[0] VDD VSS VSS RDWL S55NLLGSPH_X512Y16D32_BITCELL_RDWL2B
XI2 NET44[0] NET47[0] VDD VSS RDWL VSS S55NLLGSPH_X512Y16D32_BITCELL_RDWL2B
XI3 NET44[1] NET47[1] VDD VSS RDWL VSS S55NLLGSPH_X512Y16D32_BITCELL_RDWL2B
XI4 NET47[0] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI5 NET47[1] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI6 BL[1] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI7 BL[0] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI8 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI9 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[3] WL[2] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI10 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[5] WL[4] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI11 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[7] WL[6] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI12 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[9] WL[8] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI13 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[11] WL[10] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI14 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[13] WL[12] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI15 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[15] WL[14] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI16 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[17] WL[16] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI17 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[19] WL[18] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI18 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[21] WL[20] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI19 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[23] WL[22] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI20 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[25] WL[24] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI21 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[27] WL[26] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI22 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[29] WL[28] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI23 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[31] WL[30] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI24 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[33] WL[32] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI25 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[35] WL[34] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI26 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[37] WL[36] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI27 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[39] WL[38] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI28 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[41] WL[40] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI29 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[43] WL[42] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI30 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[45] WL[44] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI31 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[47] WL[46] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI32 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[49] WL[48] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI33 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[51] WL[50] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI34 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[53] WL[52] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI35 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[55] WL[54] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI36 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[57] WL[56] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI37 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[59] WL[58] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI38 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[61] WL[60] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI39 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[63] WL[62] S55NLLGSPH_X512Y16D32_BITCELL2X2
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN BL[1] BL[0] BLX[1] BLX[0] RDWL RWL[0] RWL[1] VDD VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0]
XI0 BL[1] BL[0] BLX[1] BLX[0] RWL[0] RWL[1] VDD VSS WL[63] WL[62]
+WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52]
+WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42]
+WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32]
+WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22]
+WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12]
+WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2]
+WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL66X2A_RED
XI1 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[127] WL[126] WL[125] WL[124]
+WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114]
+WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104]
+WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94]
+WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84]
+WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74]
+WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] S55NLLGSPH_X512Y16D32_BITCELL64X2B
XI2 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[191] WL[190] WL[189] WL[188]
+WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178]
+WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168]
+WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158]
+WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148]
+WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138]
+WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] S55NLLGSPH_X512Y16D32_BITCELL64X2A
XI3 BL[1] BL[0] BLX[1] BLX[0] RDWL VDD VSS WL[255] WL[254] WL[253]
+WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243]
+WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223]
+WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213]
+WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203]
+WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] S55NLLGSPH_X512Y16D32_BITCELL68X2B_TOP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_UP
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_UP BL[1] BL[0] BLX[1] BLX[0] RWL[0] RWL[1] VDD VSS WL[255] WL[254]
+WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244]
+WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234]
+WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224]
+WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214]
+WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204]
+WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194]
+WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184]
+WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174]
+WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164]
+WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154]
+WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144]
+WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134]
+WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124]
+WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114]
+WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104]
+WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94]
+WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84]
+WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74]
+WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64]
+WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54]
+WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44]
+WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34]
+WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24]
+WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14]
+WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4]
+WL[3] WL[2] WL[1] WL[0]
XI0 BL[1] BL[0] BLX[1] BLX[0] RWL[0] RWL[1] VDD VSS WL[63] WL[62]
+WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52]
+WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42]
+WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32]
+WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22]
+WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12]
+WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2]
+WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL66X2A_RED
XI1 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[127] WL[126] WL[125] WL[124]
+WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114]
+WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104]
+WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94]
+WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84]
+WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74]
+WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] S55NLLGSPH_X512Y16D32_BITCELL64X2B
XI2 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[191] WL[190] WL[189] WL[188]
+WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178]
+WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168]
+WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158]
+WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148]
+WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138]
+WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] S55NLLGSPH_X512Y16D32_BITCELL64X2A
XI3 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[255] WL[254] WL[253] WL[252]
+WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243] WL[242]
+WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233] WL[232]
+WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223] WL[222]
+WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213] WL[212]
+WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] WL[202]
+WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] S55NLLGSPH_X512Y16D32_BITCELL64X2B
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_YMX16SAWR
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_YMX16SAWR CLK CLKX DATA DOUT LBL[15] LBL[14] LBL[13] LBL[12] LBL[11] LBL[10]
+LBL[9] LBL[8] LBL[7] LBL[6] LBL[5] LBL[4] LBL[3] LBL[2] LBL[1] LBL[0]
+LBLX[15] LBLX[14] LBLX[13] LBLX[12] LBLX[11] LBLX[10] LBLX[9] LBLX[8] LBLX[7] LBLX[6]
+LBLX[5] LBLX[4] LBLX[3] LBLX[2] LBLX[1] LBLX[0] SACK1 SACK4 UBL[15] UBL[14]
+UBL[13] UBL[12] UBL[11] UBL[10] UBL[9] UBL[8] UBL[7] UBL[6] UBL[5] UBL[4]
+UBL[3] UBL[2] UBL[1] UBL[0] UBLX[15] UBLX[14] UBLX[13] UBLX[12] UBLX[11] UBLX[10]
+UBLX[9] UBLX[8] UBLX[7] UBLX[6] UBLX[5] UBLX[4] UBLX[3] UBLX[2] UBLX[1] UBLX[0]
+VDD VSS WE YAX YX[7] YX[6] YX[5] YX[4] YX[3] YX[2]
+YX[1] YX[0] ZAS ZASX
M0 LBL[0] 199 11 VSS N12LL L=6E-08 W=7.5E-07 $X=205 $Y=3205 $D=0
M1 11 199 LBL[0] VSS N12LL L=6E-08 W=7.5E-07 $X=205 $Y=3485 $D=0
M2 LBLX[0] 169 11 VSS N12LL L=6E-08 W=7.5E-07 $X=205 $Y=3765 $D=0
M3 11 169 LBLX[0] VSS N12LL L=6E-08 W=7.5E-07 $X=205 $Y=4045 $D=0
M4 UBLX[0] 169 12 VSS N12LL L=6E-08 W=7.5E-07 $X=205 $Y=29590 $D=0
M5 12 169 UBLX[0] VSS N12LL L=6E-08 W=7.5E-07 $X=205 $Y=29870 $D=0
M6 UBL[0] 199 12 VSS N12LL L=6E-08 W=7.5E-07 $X=205 $Y=30150 $D=0
M7 12 199 UBL[0] VSS N12LL L=6E-08 W=7.5E-07 $X=205 $Y=30430 $D=0
M8 VSS 14 1 VSS N12LL L=6E-08 W=8E-07 $X=250 $Y=9435 $D=0
M9 VSS 15 2 VSS N12LL L=6E-08 W=8E-07 $X=250 $Y=23460 $D=0
M10 VSS 1 11 VSS N12LL L=6E-08 W=1.5E-06 $X=310 $Y=4995 $D=0
M11 19 31 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=310 $Y=5265 $D=0
M12 VSS 32 20 VSS N12LL L=6E-08 W=1.5E-06 $X=310 $Y=28370 $D=0
M13 12 2 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=310 $Y=28640 $D=0
M14 16 YX[0] VSS VSS N12LL L=6E-08 W=6E-07 $X=320 $Y=22585 $D=0
M15 276 9 VSS VSS N12LL L=6E-08 W=8E-07 $X=530 $Y=9435 $D=0
M16 277 10 VSS VSS N12LL L=6E-08 W=8E-07 $X=530 $Y=23460 $D=0
M17 14 16 276 VSS N12LL L=6E-08 W=8E-07 $X=720 $Y=9435 $D=0
M18 15 16 277 VSS N12LL L=6E-08 W=8E-07 $X=720 $Y=23460 $D=0
M19 LBL[1] 199 19 VSS N12LL L=6E-08 W=7.5E-07 $X=1145 $Y=3205 $D=0
M20 19 199 LBL[1] VSS N12LL L=6E-08 W=7.5E-07 $X=1145 $Y=3485 $D=0
M21 LBLX[1] 169 19 VSS N12LL L=6E-08 W=7.5E-07 $X=1145 $Y=3765 $D=0
M22 19 169 LBLX[1] VSS N12LL L=6E-08 W=7.5E-07 $X=1145 $Y=4045 $D=0
M23 UBLX[1] 169 20 VSS N12LL L=6E-08 W=7.5E-07 $X=1145 $Y=29590 $D=0
M24 20 169 UBLX[1] VSS N12LL L=6E-08 W=7.5E-07 $X=1145 $Y=29870 $D=0
M25 UBL[1] 199 20 VSS N12LL L=6E-08 W=7.5E-07 $X=1145 $Y=30150 $D=0
M26 20 199 UBL[1] VSS N12LL L=6E-08 W=7.5E-07 $X=1145 $Y=30430 $D=0
M27 VSS YAX 17 VSS N12LL L=6E-08 W=4E-07 $X=1240 $Y=14940 $D=0
M28 VSS YAX 18 VSS N12LL L=6E-08 W=4E-07 $X=1240 $Y=19365 $D=0
M29 279 16 29 VSS N12LL L=6E-08 W=8E-07 $X=1320 $Y=9435 $D=0
M30 280 16 30 VSS N12LL L=6E-08 W=8E-07 $X=1320 $Y=23460 $D=0
M31 VSS 26 279 VSS N12LL L=6E-08 W=8E-07 $X=1510 $Y=9435 $D=0
M32 VSS 27 280 VSS N12LL L=6E-08 W=8E-07 $X=1510 $Y=23460 $D=0
M33 9 35 VSS VSS N12LL L=6E-08 W=4E-07 $X=1530 $Y=14940 $D=0
M34 10 39 VSS VSS N12LL L=6E-08 W=4E-07 $X=1530 $Y=19365 $D=0
M35 31 29 VSS VSS N12LL L=6E-08 W=8E-07 $X=1790 $Y=9435 $D=0
M36 32 30 VSS VSS N12LL L=6E-08 W=8E-07 $X=1790 $Y=23460 $D=0
M37 VSS 17 9 VSS N12LL L=6E-08 W=4E-07 $X=1820 $Y=14940 $D=0
M38 VSS 18 10 VSS N12LL L=6E-08 W=4E-07 $X=1820 $Y=19365 $D=0
M39 9 17 VSS VSS N12LL L=6E-08 W=4E-07 $X=2110 $Y=14940 $D=0
M40 10 18 VSS VSS N12LL L=6E-08 W=4E-07 $X=2110 $Y=19365 $D=0
M41 VSS ZAS 36 VSS N12LL L=6E-08 W=4E-07 $X=2135 $Y=16070 $D=0
M42 LBL[3] 199 42 VSS N12LL L=6E-08 W=7.5E-07 $X=2305 $Y=3205 $D=0
M43 42 199 LBL[3] VSS N12LL L=6E-08 W=7.5E-07 $X=2305 $Y=3485 $D=0
M44 LBLX[3] 169 42 VSS N12LL L=6E-08 W=7.5E-07 $X=2305 $Y=3765 $D=0
M45 42 169 LBLX[3] VSS N12LL L=6E-08 W=7.5E-07 $X=2305 $Y=4045 $D=0
M46 UBLX[3] 169 43 VSS N12LL L=6E-08 W=7.5E-07 $X=2305 $Y=29590 $D=0
M47 43 169 UBLX[3] VSS N12LL L=6E-08 W=7.5E-07 $X=2305 $Y=29870 $D=0
M48 UBL[3] 199 43 VSS N12LL L=6E-08 W=7.5E-07 $X=2305 $Y=30150 $D=0
M49 43 199 UBL[3] VSS N12LL L=6E-08 W=7.5E-07 $X=2305 $Y=30430 $D=0
M50 VSS 45 33 VSS N12LL L=6E-08 W=8E-07 $X=2350 $Y=9435 $D=0
M51 VSS 46 34 VSS N12LL L=6E-08 W=8E-07 $X=2350 $Y=23460 $D=0
M52 VSS 58 47 VSS N12LL L=6E-08 W=1.5E-06 $X=2390 $Y=4995 $D=0
M53 42 33 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=2390 $Y=5265 $D=0
M54 VSS 34 43 VSS N12LL L=6E-08 W=1.5E-06 $X=2390 $Y=28370 $D=0
M55 48 59 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=2390 $Y=28640 $D=0
M56 VSS 35 9 VSS N12LL L=6E-08 W=4E-07 $X=2400 $Y=14940 $D=0
M57 VSS 39 10 VSS N12LL L=6E-08 W=4E-07 $X=2400 $Y=19365 $D=0
M58 35 36 VSS VSS N12LL L=6E-08 W=4E-07 $X=2455 $Y=16070 $D=0
M59 281 26 VSS VSS N12LL L=6E-08 W=8E-07 $X=2630 $Y=9435 $D=0
M60 282 27 VSS VSS N12LL L=6E-08 W=8E-07 $X=2630 $Y=23460 $D=0
M61 9 35 VSS VSS N12LL L=6E-08 W=4E-07 $X=2690 $Y=14940 $D=0
M62 10 39 VSS VSS N12LL L=6E-08 W=4E-07 $X=2690 $Y=19365 $D=0
M63 VSS 36 35 VSS N12LL L=6E-08 W=4E-07 $X=2725 $Y=16070 $D=0
M64 45 44 281 VSS N12LL L=6E-08 W=8E-07 $X=2820 $Y=9435 $D=0
M65 46 44 282 VSS N12LL L=6E-08 W=8E-07 $X=2820 $Y=23460 $D=0
M66 VSS 17 9 VSS N12LL L=6E-08 W=4E-07 $X=2980 $Y=14940 $D=0
M67 VSS 18 10 VSS N12LL L=6E-08 W=4E-07 $X=2980 $Y=19365 $D=0
M68 39 55 VSS VSS N12LL L=6E-08 W=4E-07 $X=2995 $Y=16070 $D=0
M69 LBL[2] 199 47 VSS N12LL L=6E-08 W=7.5E-07 $X=3245 $Y=3205 $D=0
M70 47 199 LBL[2] VSS N12LL L=6E-08 W=7.5E-07 $X=3245 $Y=3485 $D=0
M71 LBLX[2] 169 47 VSS N12LL L=6E-08 W=7.5E-07 $X=3245 $Y=3765 $D=0
M72 47 169 LBLX[2] VSS N12LL L=6E-08 W=7.5E-07 $X=3245 $Y=4045 $D=0
M73 UBLX[2] 169 48 VSS N12LL L=6E-08 W=7.5E-07 $X=3245 $Y=29590 $D=0
M74 48 169 UBLX[2] VSS N12LL L=6E-08 W=7.5E-07 $X=3245 $Y=29870 $D=0
M75 UBL[2] 199 48 VSS N12LL L=6E-08 W=7.5E-07 $X=3245 $Y=30150 $D=0
M76 48 199 UBL[2] VSS N12LL L=6E-08 W=7.5E-07 $X=3245 $Y=30430 $D=0
M77 VSS 55 39 VSS N12LL L=6E-08 W=4E-07 $X=3265 $Y=16070 $D=0
M78 9 17 VSS VSS N12LL L=6E-08 W=4E-07 $X=3270 $Y=14940 $D=0
M79 10 18 VSS VSS N12LL L=6E-08 W=4E-07 $X=3270 $Y=19365 $D=0
M80 44 YX[1] VSS VSS N12LL L=6E-08 W=6E-07 $X=3280 $Y=22585 $D=0
M81 283 44 56 VSS N12LL L=6E-08 W=8E-07 $X=3420 $Y=9435 $D=0
M82 284 44 57 VSS N12LL L=6E-08 W=8E-07 $X=3420 $Y=23460 $D=0
M83 VSS 35 9 VSS N12LL L=6E-08 W=4E-07 $X=3560 $Y=14940 $D=0
M84 VSS 39 10 VSS N12LL L=6E-08 W=4E-07 $X=3560 $Y=19365 $D=0
M85 55 ZASX VSS VSS N12LL L=6E-08 W=4E-07 $X=3585 $Y=16070 $D=0
M86 VSS 9 283 VSS N12LL L=6E-08 W=8E-07 $X=3610 $Y=9435 $D=0
M87 VSS 10 284 VSS N12LL L=6E-08 W=8E-07 $X=3610 $Y=23460 $D=0
M88 26 35 VSS VSS N12LL L=6E-08 W=4E-07 $X=3850 $Y=14940 $D=0
M89 27 39 VSS VSS N12LL L=6E-08 W=4E-07 $X=3850 $Y=19365 $D=0
M90 58 56 VSS VSS N12LL L=6E-08 W=8E-07 $X=3890 $Y=9435 $D=0
M91 59 57 VSS VSS N12LL L=6E-08 W=8E-07 $X=3890 $Y=23460 $D=0
M92 VSS 9 26 VSS N12LL L=6E-08 W=4E-07 $X=4140 $Y=14940 $D=0
M93 VSS 10 27 VSS N12LL L=6E-08 W=4E-07 $X=4140 $Y=19365 $D=0
M94 VSS SACK4 65 VSS N12LL L=6E-08 W=4E-07 $X=4240 $Y=16180 $D=0
M95 LBL[4] 199 68 VSS N12LL L=6E-08 W=7.5E-07 $X=4405 $Y=3205 $D=0
M96 68 199 LBL[4] VSS N12LL L=6E-08 W=7.5E-07 $X=4405 $Y=3485 $D=0
M97 LBLX[4] 169 68 VSS N12LL L=6E-08 W=7.5E-07 $X=4405 $Y=3765 $D=0
M98 68 169 LBLX[4] VSS N12LL L=6E-08 W=7.5E-07 $X=4405 $Y=4045 $D=0
M99 UBLX[4] 169 69 VSS N12LL L=6E-08 W=7.5E-07 $X=4405 $Y=29590 $D=0
M100 69 169 UBLX[4] VSS N12LL L=6E-08 W=7.5E-07 $X=4405 $Y=29870 $D=0
M101 UBL[4] 199 69 VSS N12LL L=6E-08 W=7.5E-07 $X=4405 $Y=30150 $D=0
M102 69 199 UBL[4] VSS N12LL L=6E-08 W=7.5E-07 $X=4405 $Y=30430 $D=0
M103 26 9 VSS VSS N12LL L=6E-08 W=4E-07 $X=4430 $Y=14940 $D=0
M104 27 10 VSS VSS N12LL L=6E-08 W=4E-07 $X=4430 $Y=19365 $D=0
M105 VSS 70 61 VSS N12LL L=6E-08 W=8E-07 $X=4450 $Y=9435 $D=0
M106 VSS 71 62 VSS N12LL L=6E-08 W=8E-07 $X=4450 $Y=23460 $D=0
M107 VSS 61 68 VSS N12LL L=6E-08 W=1.5E-06 $X=4510 $Y=4995 $D=0
M108 74 82 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=4510 $Y=5265 $D=0
M109 VSS 83 75 VSS N12LL L=6E-08 W=1.5E-06 $X=4510 $Y=28370 $D=0
M110 69 62 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=4510 $Y=28640 $D=0
M111 72 YX[2] VSS VSS N12LL L=6E-08 W=6E-07 $X=4520 $Y=22585 $D=0
M112 102 65 VSS VSS N12LL L=6E-08 W=4E-07 $X=4540 $Y=16180 $D=0
M113 VSS 35 26 VSS N12LL L=6E-08 W=4E-07 $X=4720 $Y=14940 $D=0
M114 VSS 39 27 VSS N12LL L=6E-08 W=4E-07 $X=4720 $Y=19365 $D=0
M115 285 9 VSS VSS N12LL L=6E-08 W=8E-07 $X=4730 $Y=9435 $D=0
M116 286 10 VSS VSS N12LL L=6E-08 W=8E-07 $X=4730 $Y=23460 $D=0
M117 VSS 65 102 VSS N12LL L=6E-08 W=4E-07 $X=4840 $Y=16180 $D=0
M118 70 72 285 VSS N12LL L=6E-08 W=8E-07 $X=4920 $Y=9435 $D=0
M119 71 72 286 VSS N12LL L=6E-08 W=8E-07 $X=4920 $Y=23460 $D=0
M120 26 35 VSS VSS N12LL L=6E-08 W=4E-07 $X=5010 $Y=14940 $D=0
M121 27 39 VSS VSS N12LL L=6E-08 W=4E-07 $X=5010 $Y=19365 $D=0
M122 VSS 9 26 VSS N12LL L=6E-08 W=4E-07 $X=5300 $Y=14940 $D=0
M123 VSS 10 27 VSS N12LL L=6E-08 W=4E-07 $X=5300 $Y=19365 $D=0
M124 LBL[5] 199 74 VSS N12LL L=6E-08 W=7.5E-07 $X=5345 $Y=3205 $D=0
M125 74 199 LBL[5] VSS N12LL L=6E-08 W=7.5E-07 $X=5345 $Y=3485 $D=0
M126 LBLX[5] 169 74 VSS N12LL L=6E-08 W=7.5E-07 $X=5345 $Y=3765 $D=0
M127 74 169 LBLX[5] VSS N12LL L=6E-08 W=7.5E-07 $X=5345 $Y=4045 $D=0
M128 UBLX[5] 169 75 VSS N12LL L=6E-08 W=7.5E-07 $X=5345 $Y=29590 $D=0
M129 75 169 UBLX[5] VSS N12LL L=6E-08 W=7.5E-07 $X=5345 $Y=29870 $D=0
M130 UBL[5] 199 75 VSS N12LL L=6E-08 W=7.5E-07 $X=5345 $Y=30150 $D=0
M131 75 199 UBL[5] VSS N12LL L=6E-08 W=7.5E-07 $X=5345 $Y=30430 $D=0
M132 287 72 80 VSS N12LL L=6E-08 W=8E-07 $X=5520 $Y=9435 $D=0
M133 288 72 81 VSS N12LL L=6E-08 W=8E-07 $X=5520 $Y=23460 $D=0
M134 VSS 26 287 VSS N12LL L=6E-08 W=8E-07 $X=5710 $Y=9435 $D=0
M135 VSS 27 288 VSS N12LL L=6E-08 W=8E-07 $X=5710 $Y=23460 $D=0
M136 82 80 VSS VSS N12LL L=6E-08 W=8E-07 $X=5990 $Y=9435 $D=0
M137 83 81 VSS VSS N12LL L=6E-08 W=8E-07 $X=5990 $Y=23460 $D=0
M138 LBL[7] 199 90 VSS N12LL L=6E-08 W=7.5E-07 $X=6505 $Y=3205 $D=0
M139 90 199 LBL[7] VSS N12LL L=6E-08 W=7.5E-07 $X=6505 $Y=3485 $D=0
M140 LBLX[7] 169 90 VSS N12LL L=6E-08 W=7.5E-07 $X=6505 $Y=3765 $D=0
M141 90 169 LBLX[7] VSS N12LL L=6E-08 W=7.5E-07 $X=6505 $Y=4045 $D=0
M142 UBLX[7] 169 91 VSS N12LL L=6E-08 W=7.5E-07 $X=6505 $Y=29590 $D=0
M143 91 169 UBLX[7] VSS N12LL L=6E-08 W=7.5E-07 $X=6505 $Y=29870 $D=0
M144 UBL[7] 199 91 VSS N12LL L=6E-08 W=7.5E-07 $X=6505 $Y=30150 $D=0
M145 91 199 UBL[7] VSS N12LL L=6E-08 W=7.5E-07 $X=6505 $Y=30430 $D=0
M146 VSS 92 84 VSS N12LL L=6E-08 W=8E-07 $X=6550 $Y=9435 $D=0
M147 VSS 93 85 VSS N12LL L=6E-08 W=8E-07 $X=6550 $Y=23460 $D=0
M148 VSS 111 DOUT VSS N12LL L=6E-08 W=5E-07 $X=6585 $Y=15025 $D=0
M149 VSS 107 96 VSS N12LL L=6E-08 W=1.5E-06 $X=6590 $Y=4995 $D=0
M150 90 84 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=6590 $Y=5265 $D=0
M151 VSS 85 91 VSS N12LL L=6E-08 W=1.5E-06 $X=6590 $Y=28370 $D=0
M152 97 108 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=6590 $Y=28640 $D=0
M153 289 26 VSS VSS N12LL L=6E-08 W=8E-07 $X=6830 $Y=9435 $D=0
M154 290 27 VSS VSS N12LL L=6E-08 W=8E-07 $X=6830 $Y=23460 $D=0
M155 DOUT 111 VSS VSS N12LL L=6E-08 W=5E-07 $X=6875 $Y=15025 $D=0
M156 92 94 289 VSS N12LL L=6E-08 W=8E-07 $X=7020 $Y=9435 $D=0
M157 93 94 290 VSS N12LL L=6E-08 W=8E-07 $X=7020 $Y=23460 $D=0
M158 103 116 133 VSS N12LL L=1E-07 W=7.55E-07 $X=7055 $Y=17005 $D=0
M159 VSS 111 DOUT VSS N12LL L=6E-08 W=5E-07 $X=7165 $Y=15025 $D=0
M160 133 116 103 VSS N12LL L=1E-07 W=7.55E-07 $X=7425 $Y=17005 $D=0
M161 LBL[6] 199 96 VSS N12LL L=6E-08 W=7.5E-07 $X=7445 $Y=3205 $D=0
M162 96 199 LBL[6] VSS N12LL L=6E-08 W=7.5E-07 $X=7445 $Y=3485 $D=0
M163 LBLX[6] 169 96 VSS N12LL L=6E-08 W=7.5E-07 $X=7445 $Y=3765 $D=0
M164 96 169 LBLX[6] VSS N12LL L=6E-08 W=7.5E-07 $X=7445 $Y=4045 $D=0
M165 UBLX[6] 169 97 VSS N12LL L=6E-08 W=7.5E-07 $X=7445 $Y=29590 $D=0
M166 97 169 UBLX[6] VSS N12LL L=6E-08 W=7.5E-07 $X=7445 $Y=29870 $D=0
M167 UBL[6] 199 97 VSS N12LL L=6E-08 W=7.5E-07 $X=7445 $Y=30150 $D=0
M168 97 199 UBL[6] VSS N12LL L=6E-08 W=7.5E-07 $X=7445 $Y=30430 $D=0
M169 94 YX[3] VSS VSS N12LL L=6E-08 W=6E-07 $X=7480 $Y=22585 $D=0
M170 291 94 105 VSS N12LL L=6E-08 W=8E-07 $X=7620 $Y=9435 $D=0
M171 292 94 106 VSS N12LL L=6E-08 W=8E-07 $X=7620 $Y=23460 $D=0
M172 103 116 133 VSS N12LL L=1E-07 W=7.55E-07 $X=7795 $Y=17005 $D=0
M173 VSS 9 291 VSS N12LL L=6E-08 W=8E-07 $X=7810 $Y=9435 $D=0
M174 VSS 10 292 VSS N12LL L=6E-08 W=8E-07 $X=7810 $Y=23460 $D=0
M175 293 102 VSS VSS N12LL L=6E-08 W=1E-06 $X=7900 $Y=16325 $D=0
M176 133 139 293 VSS N12LL L=6E-08 W=1E-06 $X=7900 $Y=16535 $D=0
M177 294 103 111 VSS N12LL L=6E-08 W=1E-06 $X=7930 $Y=14925 $D=0
M178 107 105 VSS VSS N12LL L=6E-08 W=8E-07 $X=8090 $Y=9435 $D=0
M179 108 106 VSS VSS N12LL L=6E-08 W=8E-07 $X=8090 $Y=23460 $D=0
M180 133 116 103 VSS N12LL L=1E-07 W=7.55E-07 $X=8165 $Y=17005 $D=0
M181 VSS 121 294 VSS N12LL L=6E-08 W=1E-06 $X=8220 $Y=14925 $D=0
M182 295 111 VSS VSS N12LL L=6E-08 W=1E-06 $X=8510 $Y=14925 $D=0
M183 116 103 133 VSS N12LL L=1E-07 W=7.55E-07 $X=8535 $Y=17005 $D=0
M184 LBL[8] 199 119 VSS N12LL L=6E-08 W=7.5E-07 $X=8605 $Y=3205 $D=0
M185 119 199 LBL[8] VSS N12LL L=6E-08 W=7.5E-07 $X=8605 $Y=3485 $D=0
M186 LBLX[8] 169 119 VSS N12LL L=6E-08 W=7.5E-07 $X=8605 $Y=3765 $D=0
M187 119 169 LBLX[8] VSS N12LL L=6E-08 W=7.5E-07 $X=8605 $Y=4045 $D=0
M188 UBLX[8] 169 120 VSS N12LL L=6E-08 W=7.5E-07 $X=8605 $Y=29590 $D=0
M189 120 169 UBLX[8] VSS N12LL L=6E-08 W=7.5E-07 $X=8605 $Y=29870 $D=0
M190 UBL[8] 199 120 VSS N12LL L=6E-08 W=7.5E-07 $X=8605 $Y=30150 $D=0
M191 120 199 UBL[8] VSS N12LL L=6E-08 W=7.5E-07 $X=8605 $Y=30430 $D=0
M192 VSS 124 112 VSS N12LL L=6E-08 W=8E-07 $X=8650 $Y=9435 $D=0
M193 VSS 125 113 VSS N12LL L=6E-08 W=8E-07 $X=8650 $Y=23460 $D=0
M194 VSS 112 119 VSS N12LL L=6E-08 W=1.5E-06 $X=8710 $Y=4995 $D=0
M195 127 137 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=8710 $Y=5265 $D=0
M196 VSS 138 128 VSS N12LL L=6E-08 W=1.5E-06 $X=8710 $Y=28370 $D=0
M197 120 113 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=8710 $Y=28640 $D=0
M198 VSS YX[4] 126 VSS N12LL L=6E-08 W=6E-07 $X=8720 $Y=11050 $D=0
M199 121 116 295 VSS N12LL L=6E-08 W=1E-06 $X=8800 $Y=14925 $D=0
M200 133 103 116 VSS N12LL L=1E-07 W=7.55E-07 $X=8905 $Y=17005 $D=0
M201 297 9 VSS VSS N12LL L=6E-08 W=8E-07 $X=8930 $Y=9435 $D=0
M202 298 10 VSS VSS N12LL L=6E-08 W=8E-07 $X=8930 $Y=23460 $D=0
M203 124 126 297 VSS N12LL L=6E-08 W=8E-07 $X=9120 $Y=9435 $D=0
M204 125 126 298 VSS N12LL L=6E-08 W=8E-07 $X=9120 $Y=23460 $D=0
M205 116 103 133 VSS N12LL L=1E-07 W=7.55E-07 $X=9275 $Y=17005 $D=0
M206 LBL[9] 199 127 VSS N12LL L=6E-08 W=7.5E-07 $X=9545 $Y=3205 $D=0
M207 127 199 LBL[9] VSS N12LL L=6E-08 W=7.5E-07 $X=9545 $Y=3485 $D=0
M208 LBLX[9] 169 127 VSS N12LL L=6E-08 W=7.5E-07 $X=9545 $Y=3765 $D=0
M209 127 169 LBLX[9] VSS N12LL L=6E-08 W=7.5E-07 $X=9545 $Y=4045 $D=0
M210 UBLX[9] 169 128 VSS N12LL L=6E-08 W=7.5E-07 $X=9545 $Y=29590 $D=0
M211 128 169 UBLX[9] VSS N12LL L=6E-08 W=7.5E-07 $X=9545 $Y=29870 $D=0
M212 UBL[9] 199 128 VSS N12LL L=6E-08 W=7.5E-07 $X=9545 $Y=30150 $D=0
M213 128 199 UBL[9] VSS N12LL L=6E-08 W=7.5E-07 $X=9545 $Y=30430 $D=0
M214 133 103 116 VSS N12LL L=1E-07 W=7.55E-07 $X=9645 $Y=17005 $D=0
M215 299 126 134 VSS N12LL L=6E-08 W=8E-07 $X=9720 $Y=9435 $D=0
M216 300 126 135 VSS N12LL L=6E-08 W=8E-07 $X=9720 $Y=23460 $D=0
M217 VSS 26 299 VSS N12LL L=6E-08 W=8E-07 $X=9910 $Y=9435 $D=0
M218 VSS 27 300 VSS N12LL L=6E-08 W=8E-07 $X=9910 $Y=23460 $D=0
M219 VSS VSS DATA VSS N12LL L=6E-08 W=2E-07 $X=9980 $Y=15575 $D=0
M220 137 134 VSS VSS N12LL L=6E-08 W=8E-07 $X=10190 $Y=9435 $D=0
M221 138 135 VSS VSS N12LL L=6E-08 W=8E-07 $X=10190 $Y=23460 $D=0
M222 VSS DATA 140 VSS N12LL L=6E-08 W=4E-07 $X=10195 $Y=14885 $D=0
M223 150 140 VSS VSS N12LL L=3E-07 W=4E-07 $X=10545 $Y=14885 $D=0
M224 VSS 147 139 VSS N12LL L=6E-08 W=5E-07 $X=10590 $Y=19250 $D=0
M225 LBL[11] 199 148 VSS N12LL L=6E-08 W=7.5E-07 $X=10705 $Y=3205 $D=0
M226 148 199 LBL[11] VSS N12LL L=6E-08 W=7.5E-07 $X=10705 $Y=3485 $D=0
M227 LBLX[11] 169 148 VSS N12LL L=6E-08 W=7.5E-07 $X=10705 $Y=3765 $D=0
M228 148 169 LBLX[11] VSS N12LL L=6E-08 W=7.5E-07 $X=10705 $Y=4045 $D=0
M229 UBLX[11] 169 149 VSS N12LL L=6E-08 W=7.5E-07 $X=10705 $Y=29590 $D=0
M230 149 169 UBLX[11] VSS N12LL L=6E-08 W=7.5E-07 $X=10705 $Y=29870 $D=0
M231 UBL[11] 199 149 VSS N12LL L=6E-08 W=7.5E-07 $X=10705 $Y=30150 $D=0
M232 149 199 UBL[11] VSS N12LL L=6E-08 W=7.5E-07 $X=10705 $Y=30430 $D=0
M233 VSS 151 141 VSS N12LL L=6E-08 W=8E-07 $X=10750 $Y=9435 $D=0
M234 VSS 152 142 VSS N12LL L=6E-08 W=8E-07 $X=10750 $Y=23460 $D=0
M235 VSS 166 154 VSS N12LL L=6E-08 W=1.5E-06 $X=10790 $Y=4995 $D=0
M236 148 141 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=10790 $Y=5265 $D=0
M237 VSS 142 149 VSS N12LL L=6E-08 W=1.5E-06 $X=10790 $Y=28370 $D=0
M238 155 167 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=10790 $Y=28640 $D=0
M239 147 SACK1 VSS VSS N12LL L=6E-08 W=4E-07 $X=10890 $Y=19350 $D=0
M240 301 26 VSS VSS N12LL L=6E-08 W=8E-07 $X=11030 $Y=9435 $D=0
M241 302 27 VSS VSS N12LL L=6E-08 W=8E-07 $X=11030 $Y=23460 $D=0
M242 151 153 301 VSS N12LL L=6E-08 W=8E-07 $X=11220 $Y=9435 $D=0
M243 152 153 302 VSS N12LL L=6E-08 W=8E-07 $X=11220 $Y=23460 $D=0
M244 VSS 202 185 VSS N12LL L=6E-08 W=4E-07 $X=11405 $Y=16275 $D=0
M245 VSS 150 159 VSS N12LL L=2E-07 W=4E-07 $X=11505 $Y=14885 $D=0
M246 VSS 165 109 VSS N12LL L=6E-08 W=5E-07 $X=11515 $Y=19250 $D=0
M247 LBL[10] 199 154 VSS N12LL L=6E-08 W=7.5E-07 $X=11645 $Y=3205 $D=0
M248 154 199 LBL[10] VSS N12LL L=6E-08 W=7.5E-07 $X=11645 $Y=3485 $D=0
M249 LBLX[10] 169 154 VSS N12LL L=6E-08 W=7.5E-07 $X=11645 $Y=3765 $D=0
M250 154 169 LBLX[10] VSS N12LL L=6E-08 W=7.5E-07 $X=11645 $Y=4045 $D=0
M251 UBLX[10] 169 155 VSS N12LL L=6E-08 W=7.5E-07 $X=11645 $Y=29590 $D=0
M252 155 169 UBLX[10] VSS N12LL L=6E-08 W=7.5E-07 $X=11645 $Y=29870 $D=0
M253 UBL[10] 199 155 VSS N12LL L=6E-08 W=7.5E-07 $X=11645 $Y=30150 $D=0
M254 155 199 UBL[10] VSS N12LL L=6E-08 W=7.5E-07 $X=11645 $Y=30430 $D=0
M255 VSS YX[5] 153 VSS N12LL L=6E-08 W=6E-07 $X=11680 $Y=11050 $D=0
M256 304 SACK1 VSS VSS N12LL L=6E-08 W=4E-07 $X=11815 $Y=19350 $D=0
M257 305 153 163 VSS N12LL L=6E-08 W=8E-07 $X=11820 $Y=9435 $D=0
M258 306 153 164 VSS N12LL L=6E-08 W=8E-07 $X=11820 $Y=23460 $D=0
M259 168 159 VSS VSS N12LL L=6E-08 W=7E-07 $X=11995 $Y=14885 $D=0
M260 VSS 9 305 VSS N12LL L=6E-08 W=8E-07 $X=12010 $Y=9435 $D=0
M261 VSS 10 306 VSS N12LL L=6E-08 W=8E-07 $X=12010 $Y=23460 $D=0
M262 165 SACK4 304 VSS N12LL L=6E-08 W=4E-07 $X=12105 $Y=19350 $D=0
M263 VSS 202 172 VSS N12LL L=6E-07 W=1.2E-07 $X=12155 $Y=16555 $D=0
M264 166 163 VSS VSS N12LL L=6E-08 W=8E-07 $X=12290 $Y=9435 $D=0
M265 167 164 VSS VSS N12LL L=6E-08 W=8E-07 $X=12290 $Y=23460 $D=0
M266 172 CLKX 168 VSS N12LL L=6E-08 W=7E-07 $X=12675 $Y=14885 $D=0
M267 LBL[12] 199 179 VSS N12LL L=6E-08 W=7.5E-07 $X=12805 $Y=3205 $D=0
M268 179 199 LBL[12] VSS N12LL L=6E-08 W=7.5E-07 $X=12805 $Y=3485 $D=0
M269 LBLX[12] 169 179 VSS N12LL L=6E-08 W=7.5E-07 $X=12805 $Y=3765 $D=0
M270 179 169 LBLX[12] VSS N12LL L=6E-08 W=7.5E-07 $X=12805 $Y=4045 $D=0
M271 UBLX[12] 169 180 VSS N12LL L=6E-08 W=7.5E-07 $X=12805 $Y=29590 $D=0
M272 180 169 UBLX[12] VSS N12LL L=6E-08 W=7.5E-07 $X=12805 $Y=29870 $D=0
M273 UBL[12] 199 180 VSS N12LL L=6E-08 W=7.5E-07 $X=12805 $Y=30150 $D=0
M274 180 199 UBL[12] VSS N12LL L=6E-08 W=7.5E-07 $X=12805 $Y=30430 $D=0
M275 VSS 181 173 VSS N12LL L=6E-08 W=8E-07 $X=12850 $Y=9435 $D=0
M276 VSS 182 174 VSS N12LL L=6E-08 W=8E-07 $X=12850 $Y=23460 $D=0
M277 VSS 173 179 VSS N12LL L=6E-08 W=1.5E-06 $X=12910 $Y=4995 $D=0
M278 186 196 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=12910 $Y=5265 $D=0
M279 VSS 197 187 VSS N12LL L=6E-08 W=1.5E-06 $X=12910 $Y=28370 $D=0
M280 180 174 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=12910 $Y=28640 $D=0
M281 VSS YX[6] 183 VSS N12LL L=6E-08 W=6E-07 $X=12920 $Y=11050 $D=0
M282 169 193 VSS VSS N12LL L=6E-08 W=1E-06 $X=13040 $Y=18935 $D=0
M283 202 172 VSS VSS N12LL L=6E-08 W=5E-07 $X=13090 $Y=16175 $D=0
M284 308 9 VSS VSS N12LL L=6E-08 W=8E-07 $X=13130 $Y=9435 $D=0
M285 309 10 VSS VSS N12LL L=6E-08 W=8E-07 $X=13130 $Y=23460 $D=0
M286 188 CLKX 200 VSS N12LL L=6E-08 W=7E-07 $X=13295 $Y=14885 $D=0
M287 181 183 308 VSS N12LL L=6E-08 W=8E-07 $X=13320 $Y=9435 $D=0
M288 182 183 309 VSS N12LL L=6E-08 W=8E-07 $X=13320 $Y=23460 $D=0
M289 VSS 193 169 VSS N12LL L=6E-08 W=1E-06 $X=13330 $Y=18935 $D=0
M290 310 185 VSS VSS N12LL L=6E-08 W=1E-06 $X=13620 $Y=18935 $D=0
M291 LBL[13] 199 186 VSS N12LL L=6E-08 W=7.5E-07 $X=13745 $Y=3205 $D=0
M292 186 199 LBL[13] VSS N12LL L=6E-08 W=7.5E-07 $X=13745 $Y=3485 $D=0
M293 LBLX[13] 169 186 VSS N12LL L=6E-08 W=7.5E-07 $X=13745 $Y=3765 $D=0
M294 186 169 LBLX[13] VSS N12LL L=6E-08 W=7.5E-07 $X=13745 $Y=4045 $D=0
M295 UBLX[13] 169 187 VSS N12LL L=6E-08 W=7.5E-07 $X=13745 $Y=29590 $D=0
M296 187 169 UBLX[13] VSS N12LL L=6E-08 W=7.5E-07 $X=13745 $Y=29870 $D=0
M297 UBL[13] 199 187 VSS N12LL L=6E-08 W=7.5E-07 $X=13745 $Y=30150 $D=0
M298 187 199 UBL[13] VSS N12LL L=6E-08 W=7.5E-07 $X=13745 $Y=30430 $D=0
M299 VSS 200 212 VSS N12LL L=6E-08 W=4E-07 $X=13750 $Y=16275 $D=0
M300 311 183 194 VSS N12LL L=6E-08 W=8E-07 $X=13920 $Y=9435 $D=0
M301 312 183 195 VSS N12LL L=6E-08 W=8E-07 $X=13920 $Y=23460 $D=0
M302 193 227 310 VSS N12LL L=6E-08 W=1E-06 $X=13925 $Y=18935 $D=0
M303 VSS 198 188 VSS N12LL L=6E-08 W=7E-07 $X=13955 $Y=14885 $D=0
M304 VSS 26 311 VSS N12LL L=6E-08 W=8E-07 $X=14110 $Y=9435 $D=0
M305 VSS 27 312 VSS N12LL L=6E-08 W=8E-07 $X=14110 $Y=23460 $D=0
M306 200 212 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=14145 $Y=16555 $D=0
M307 198 207 VSS VSS N12LL L=2E-07 W=4E-07 $X=14305 $Y=14885 $D=0
M308 196 194 VSS VSS N12LL L=6E-08 W=8E-07 $X=14390 $Y=9435 $D=0
M309 197 195 VSS VSS N12LL L=6E-08 W=8E-07 $X=14390 $Y=23460 $D=0
M310 313 227 201 VSS N12LL L=6E-08 W=1E-06 $X=14605 $Y=18935 $D=0
M311 LBL[15] 199 210 VSS N12LL L=6E-08 W=7.5E-07 $X=14905 $Y=3205 $D=0
M312 210 199 LBL[15] VSS N12LL L=6E-08 W=7.5E-07 $X=14905 $Y=3485 $D=0
M313 LBLX[15] 169 210 VSS N12LL L=6E-08 W=7.5E-07 $X=14905 $Y=3765 $D=0
M314 210 169 LBLX[15] VSS N12LL L=6E-08 W=7.5E-07 $X=14905 $Y=4045 $D=0
M315 UBLX[15] 169 211 VSS N12LL L=6E-08 W=7.5E-07 $X=14905 $Y=29590 $D=0
M316 211 169 UBLX[15] VSS N12LL L=6E-08 W=7.5E-07 $X=14905 $Y=29870 $D=0
M317 UBL[15] 199 211 VSS N12LL L=6E-08 W=7.5E-07 $X=14905 $Y=30150 $D=0
M318 211 199 UBL[15] VSS N12LL L=6E-08 W=7.5E-07 $X=14905 $Y=30430 $D=0
M319 VSS 202 313 VSS N12LL L=6E-08 W=1E-06 $X=14910 $Y=18935 $D=0
M320 VSS 213 203 VSS N12LL L=6E-08 W=8E-07 $X=14950 $Y=9435 $D=0
M321 VSS 215 204 VSS N12LL L=6E-08 W=8E-07 $X=14950 $Y=23460 $D=0
M322 VSS 231 218 VSS N12LL L=6E-08 W=1.5E-06 $X=14990 $Y=4995 $D=0
M323 210 203 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=14990 $Y=5265 $D=0
M324 VSS 204 211 VSS N12LL L=6E-08 W=1.5E-06 $X=14990 $Y=28370 $D=0
M325 219 232 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=14990 $Y=28640 $D=0
M326 VSS 217 207 VSS N12LL L=3E-07 W=4E-07 $X=15165 $Y=14885 $D=0
M327 199 201 VSS VSS N12LL L=6E-08 W=1E-06 $X=15200 $Y=18935 $D=0
M328 314 26 VSS VSS N12LL L=6E-08 W=8E-07 $X=15230 $Y=9435 $D=0
M329 315 27 VSS VSS N12LL L=6E-08 W=8E-07 $X=15230 $Y=23460 $D=0
M330 213 214 314 VSS N12LL L=6E-08 W=8E-07 $X=15420 $Y=9435 $D=0
M331 215 214 315 VSS N12LL L=6E-08 W=8E-07 $X=15420 $Y=23460 $D=0
M332 316 212 220 VSS N12LL L=6E-08 W=4E-07 $X=15460 $Y=16125 $D=0
M333 VSS 201 199 VSS N12LL L=6E-08 W=1E-06 $X=15490 $Y=18935 $D=0
M334 217 226 VSS VSS N12LL L=6E-08 W=4E-07 $X=15755 $Y=14885 $D=0
M335 VSS WE 316 VSS N12LL L=6E-08 W=4E-07 $X=15765 $Y=16125 $D=0
M336 LBL[14] 199 218 VSS N12LL L=6E-08 W=7.5E-07 $X=15845 $Y=3205 $D=0
M337 218 199 LBL[14] VSS N12LL L=6E-08 W=7.5E-07 $X=15845 $Y=3485 $D=0
M338 LBLX[14] 169 218 VSS N12LL L=6E-08 W=7.5E-07 $X=15845 $Y=3765 $D=0
M339 218 169 LBLX[14] VSS N12LL L=6E-08 W=7.5E-07 $X=15845 $Y=4045 $D=0
M340 UBLX[14] 169 219 VSS N12LL L=6E-08 W=7.5E-07 $X=15845 $Y=29590 $D=0
M341 219 169 UBLX[14] VSS N12LL L=6E-08 W=7.5E-07 $X=15845 $Y=29870 $D=0
M342 UBL[14] 199 219 VSS N12LL L=6E-08 W=7.5E-07 $X=15845 $Y=30150 $D=0
M343 219 199 UBL[14] VSS N12LL L=6E-08 W=7.5E-07 $X=15845 $Y=30430 $D=0
M344 VSS YX[7] 214 VSS N12LL L=6E-08 W=6E-07 $X=15880 $Y=11050 $D=0
M345 318 214 228 VSS N12LL L=6E-08 W=8E-07 $X=16020 $Y=9435 $D=0
M346 319 214 229 VSS N12LL L=6E-08 W=8E-07 $X=16020 $Y=23460 $D=0
M347 227 220 VSS VSS N12LL L=6E-08 W=5E-07 $X=16055 $Y=16025 $D=0
M348 VSS 9 318 VSS N12LL L=6E-08 W=8E-07 $X=16210 $Y=9435 $D=0
M349 VSS 10 319 VSS N12LL L=6E-08 W=8E-07 $X=16210 $Y=23460 $D=0
M350 VSS 230 226 VSS N12LL L=6E-08 W=1E-06 $X=16410 $Y=14885 $D=0
M351 231 228 VSS VSS N12LL L=6E-08 W=8E-07 $X=16490 $Y=9435 $D=0
M352 232 229 VSS VSS N12LL L=6E-08 W=8E-07 $X=16490 $Y=23460 $D=0
M353 LBL[0] 1 VDD VDD P12LL L=6E-08 W=1E-06 $X=185 $Y=1635 $D=1
M354 UBL[0] 2 VDD VDD P12LL L=6E-08 W=1E-06 $X=185 $Y=31060 $D=1
M355 VDD 14 1 VDD P12LL L=6E-08 W=6E-07 $X=250 $Y=8205 $D=1
M356 VDD 15 2 VDD P12LL L=6E-08 W=6E-07 $X=250 $Y=24890 $D=1
M357 122 14 LBLX[0] VDD P12LL L=6E-08 W=6E-07 $X=295 $Y=5965 $D=1
M358 110 14 LBL[0] VDD P12LL L=6E-08 W=6E-07 $X=295 $Y=6885 $D=1
M359 110 15 UBL[0] VDD P12LL L=6E-08 W=6E-07 $X=295 $Y=26210 $D=1
M360 122 15 UBLX[0] VDD P12LL L=6E-08 W=6E-07 $X=295 $Y=27130 $D=1
M361 LBLX[0] 1 LBL[0] VDD P12LL L=6E-08 W=1E-06 $X=495 $Y=1635 $D=1
M362 UBLX[0] 2 UBL[0] VDD P12LL L=6E-08 W=1E-06 $X=495 $Y=31060 $D=1
M363 14 9 VDD VDD P12LL L=6E-08 W=6E-07 $X=530 $Y=8205 $D=1
M364 15 10 VDD VDD P12LL L=6E-08 W=6E-07 $X=530 $Y=24890 $D=1
M365 VDD 1 LBLX[0] VDD P12LL L=6E-08 W=1E-06 $X=805 $Y=1635 $D=1
M366 VDD 2 UBLX[0] VDD P12LL L=6E-08 W=1E-06 $X=805 $Y=31060 $D=1
M367 VDD 16 14 VDD P12LL L=6E-08 W=6E-07 $X=810 $Y=8205 $D=1
M368 VDD 16 15 VDD P12LL L=6E-08 W=6E-07 $X=810 $Y=24890 $D=1
M369 29 16 VDD VDD P12LL L=6E-08 W=6E-07 $X=1230 $Y=8205 $D=1
M370 30 16 VDD VDD P12LL L=6E-08 W=6E-07 $X=1230 $Y=24890 $D=1
M371 LBLX[1] 31 VDD VDD P12LL L=6E-08 W=1E-06 $X=1235 $Y=1635 $D=1
M372 UBLX[1] 32 VDD VDD P12LL L=6E-08 W=1E-06 $X=1235 $Y=31060 $D=1
M373 VDD YAX 17 VDD P12LL L=6E-08 W=8E-07 $X=1240 $Y=13360 $D=1
M374 VDD YAX 18 VDD P12LL L=6E-08 W=8E-07 $X=1240 $Y=20545 $D=1
M375 16 YX[0] VDD VDD P12LL L=6E-08 W=4E-07 $X=1380 $Y=22045 $D=1
M376 VDD YX[0] 16 VDD P12LL L=6E-08 W=4E-07 $X=1380 $Y=22315 $D=1
M377 16 YX[0] VDD VDD P12LL L=6E-08 W=4E-07 $X=1380 $Y=22585 $D=1
M378 VDD 26 29 VDD P12LL L=6E-08 W=6E-07 $X=1510 $Y=8205 $D=1
M379 VDD 27 30 VDD P12LL L=6E-08 W=6E-07 $X=1510 $Y=24890 $D=1
M380 323 35 VDD VDD P12LL L=6E-08 W=8E-07 $X=1530 $Y=13360 $D=1
M381 324 39 VDD VDD P12LL L=6E-08 W=8E-07 $X=1530 $Y=20545 $D=1
M382 LBL[1] 31 LBLX[1] VDD P12LL L=6E-08 W=1E-06 $X=1545 $Y=1635 $D=1
M383 UBL[1] 32 UBLX[1] VDD P12LL L=6E-08 W=1E-06 $X=1545 $Y=31060 $D=1
M384 LBLX[1] 29 122 VDD P12LL L=6E-08 W=6E-07 $X=1745 $Y=5965 $D=1
M385 LBL[1] 29 110 VDD P12LL L=6E-08 W=6E-07 $X=1745 $Y=6885 $D=1
M386 UBL[1] 30 110 VDD P12LL L=6E-08 W=6E-07 $X=1745 $Y=26210 $D=1
M387 UBLX[1] 30 122 VDD P12LL L=6E-08 W=6E-07 $X=1745 $Y=27130 $D=1
M388 31 29 VDD VDD P12LL L=6E-08 W=6E-07 $X=1790 $Y=8205 $D=1
M389 32 30 VDD VDD P12LL L=6E-08 W=6E-07 $X=1790 $Y=24890 $D=1
M390 9 17 323 VDD P12LL L=6E-08 W=8E-07 $X=1820 $Y=13360 $D=1
M391 10 18 324 VDD P12LL L=6E-08 W=8E-07 $X=1820 $Y=20545 $D=1
M392 VDD 31 LBL[1] VDD P12LL L=6E-08 W=1E-06 $X=1855 $Y=1635 $D=1
M393 VDD 32 UBL[1] VDD P12LL L=6E-08 W=1E-06 $X=1855 $Y=31060 $D=1
M394 325 17 9 VDD P12LL L=6E-08 W=8E-07 $X=2110 $Y=13360 $D=1
M395 326 18 10 VDD P12LL L=6E-08 W=8E-07 $X=2110 $Y=20545 $D=1
M396 VDD ZAS 36 VDD P12LL L=6E-08 W=4E-07 $X=2135 $Y=17430 $D=1
M397 LBL[3] 33 VDD VDD P12LL L=6E-08 W=1E-06 $X=2285 $Y=1635 $D=1
M398 UBL[3] 34 VDD VDD P12LL L=6E-08 W=1E-06 $X=2285 $Y=31060 $D=1
M399 VDD 45 33 VDD P12LL L=6E-08 W=6E-07 $X=2350 $Y=8205 $D=1
M400 VDD 46 34 VDD P12LL L=6E-08 W=6E-07 $X=2350 $Y=24890 $D=1
M401 122 45 LBLX[3] VDD P12LL L=6E-08 W=6E-07 $X=2395 $Y=5965 $D=1
M402 110 45 LBL[3] VDD P12LL L=6E-08 W=6E-07 $X=2395 $Y=6885 $D=1
M403 110 46 UBL[3] VDD P12LL L=6E-08 W=6E-07 $X=2395 $Y=26210 $D=1
M404 122 46 UBLX[3] VDD P12LL L=6E-08 W=6E-07 $X=2395 $Y=27130 $D=1
M405 VDD 35 325 VDD P12LL L=6E-08 W=8E-07 $X=2400 $Y=13360 $D=1
M406 VDD 39 326 VDD P12LL L=6E-08 W=8E-07 $X=2400 $Y=20545 $D=1
M407 44 YX[1] VDD VDD P12LL L=6E-08 W=4E-07 $X=2420 $Y=22045 $D=1
M408 VDD YX[1] 44 VDD P12LL L=6E-08 W=4E-07 $X=2420 $Y=22315 $D=1
M409 44 YX[1] VDD VDD P12LL L=6E-08 W=4E-07 $X=2420 $Y=22585 $D=1
M410 35 36 VDD VDD P12LL L=6E-08 W=8E-07 $X=2455 $Y=17430 $D=1
M411 LBLX[3] 33 LBL[3] VDD P12LL L=6E-08 W=1E-06 $X=2595 $Y=1635 $D=1
M412 UBLX[3] 34 UBL[3] VDD P12LL L=6E-08 W=1E-06 $X=2595 $Y=31060 $D=1
M413 45 26 VDD VDD P12LL L=6E-08 W=6E-07 $X=2630 $Y=8205 $D=1
M414 46 27 VDD VDD P12LL L=6E-08 W=6E-07 $X=2630 $Y=24890 $D=1
M415 327 35 VDD VDD P12LL L=6E-08 W=8E-07 $X=2690 $Y=13360 $D=1
M416 328 39 VDD VDD P12LL L=6E-08 W=8E-07 $X=2690 $Y=20545 $D=1
M417 VDD 36 35 VDD P12LL L=6E-08 W=8E-07 $X=2725 $Y=17430 $D=1
M418 VDD 33 LBLX[3] VDD P12LL L=6E-08 W=1E-06 $X=2905 $Y=1635 $D=1
M419 VDD 34 UBLX[3] VDD P12LL L=6E-08 W=1E-06 $X=2905 $Y=31060 $D=1
M420 VDD 44 45 VDD P12LL L=6E-08 W=6E-07 $X=2910 $Y=8205 $D=1
M421 VDD 44 46 VDD P12LL L=6E-08 W=6E-07 $X=2910 $Y=24890 $D=1
M422 9 17 327 VDD P12LL L=6E-08 W=8E-07 $X=2980 $Y=13360 $D=1
M423 10 18 328 VDD P12LL L=6E-08 W=8E-07 $X=2980 $Y=20545 $D=1
M424 39 55 VDD VDD P12LL L=6E-08 W=8E-07 $X=2995 $Y=17430 $D=1
M425 VDD 55 39 VDD P12LL L=6E-08 W=8E-07 $X=3265 $Y=17430 $D=1
M426 329 17 9 VDD P12LL L=6E-08 W=8E-07 $X=3270 $Y=13360 $D=1
M427 330 18 10 VDD P12LL L=6E-08 W=8E-07 $X=3270 $Y=20545 $D=1
M428 56 44 VDD VDD P12LL L=6E-08 W=6E-07 $X=3330 $Y=8205 $D=1
M429 57 44 VDD VDD P12LL L=6E-08 W=6E-07 $X=3330 $Y=24890 $D=1
M430 LBLX[2] 58 VDD VDD P12LL L=6E-08 W=1E-06 $X=3335 $Y=1635 $D=1
M431 UBLX[2] 59 VDD VDD P12LL L=6E-08 W=1E-06 $X=3335 $Y=31060 $D=1
M432 VDD 35 329 VDD P12LL L=6E-08 W=8E-07 $X=3560 $Y=13360 $D=1
M433 VDD 39 330 VDD P12LL L=6E-08 W=8E-07 $X=3560 $Y=20545 $D=1
M434 55 ZASX VDD VDD P12LL L=6E-08 W=4E-07 $X=3585 $Y=17430 $D=1
M435 VDD 9 56 VDD P12LL L=6E-08 W=6E-07 $X=3610 $Y=8205 $D=1
M436 VDD 10 57 VDD P12LL L=6E-08 W=6E-07 $X=3610 $Y=24890 $D=1
M437 LBL[2] 58 LBLX[2] VDD P12LL L=6E-08 W=1E-06 $X=3645 $Y=1635 $D=1
M438 UBL[2] 59 UBLX[2] VDD P12LL L=6E-08 W=1E-06 $X=3645 $Y=31060 $D=1
M439 LBLX[2] 56 122 VDD P12LL L=6E-08 W=6E-07 $X=3845 $Y=5965 $D=1
M440 LBL[2] 56 110 VDD P12LL L=6E-08 W=6E-07 $X=3845 $Y=6885 $D=1
M441 UBL[2] 57 110 VDD P12LL L=6E-08 W=6E-07 $X=3845 $Y=26210 $D=1
M442 UBLX[2] 57 122 VDD P12LL L=6E-08 W=6E-07 $X=3845 $Y=27130 $D=1
M443 331 35 VDD VDD P12LL L=6E-08 W=8E-07 $X=3850 $Y=13360 $D=1
M444 332 39 VDD VDD P12LL L=6E-08 W=8E-07 $X=3850 $Y=20545 $D=1
M445 58 56 VDD VDD P12LL L=6E-08 W=6E-07 $X=3890 $Y=8205 $D=1
M446 59 57 VDD VDD P12LL L=6E-08 W=6E-07 $X=3890 $Y=24890 $D=1
M447 VDD 58 LBL[2] VDD P12LL L=6E-08 W=1E-06 $X=3955 $Y=1635 $D=1
M448 VDD 59 UBL[2] VDD P12LL L=6E-08 W=1E-06 $X=3955 $Y=31060 $D=1
M449 26 9 331 VDD P12LL L=6E-08 W=8E-07 $X=4140 $Y=13360 $D=1
M450 27 10 332 VDD P12LL L=6E-08 W=8E-07 $X=4140 $Y=20545 $D=1
M451 VDD SACK4 65 VDD P12LL L=6E-08 W=8E-07 $X=4240 $Y=17355 $D=1
M452 LBL[4] 61 VDD VDD P12LL L=6E-08 W=1E-06 $X=4385 $Y=1635 $D=1
M453 UBL[4] 62 VDD VDD P12LL L=6E-08 W=1E-06 $X=4385 $Y=31060 $D=1
M454 333 9 26 VDD P12LL L=6E-08 W=8E-07 $X=4430 $Y=13360 $D=1
M455 334 10 27 VDD P12LL L=6E-08 W=8E-07 $X=4430 $Y=20545 $D=1
M456 VDD 70 61 VDD P12LL L=6E-08 W=6E-07 $X=4450 $Y=8205 $D=1
M457 VDD 71 62 VDD P12LL L=6E-08 W=6E-07 $X=4450 $Y=24890 $D=1
M458 122 70 LBLX[4] VDD P12LL L=6E-08 W=6E-07 $X=4495 $Y=5965 $D=1
M459 110 70 LBL[4] VDD P12LL L=6E-08 W=6E-07 $X=4495 $Y=6885 $D=1
M460 110 71 UBL[4] VDD P12LL L=6E-08 W=6E-07 $X=4495 $Y=26210 $D=1
M461 122 71 UBLX[4] VDD P12LL L=6E-08 W=6E-07 $X=4495 $Y=27130 $D=1
M462 102 65 VDD VDD P12LL L=6E-08 W=8E-07 $X=4540 $Y=17355 $D=1
M463 LBLX[4] 61 LBL[4] VDD P12LL L=6E-08 W=1E-06 $X=4695 $Y=1635 $D=1
M464 UBLX[4] 62 UBL[4] VDD P12LL L=6E-08 W=1E-06 $X=4695 $Y=31060 $D=1
M465 VDD 35 333 VDD P12LL L=6E-08 W=8E-07 $X=4720 $Y=13360 $D=1
M466 VDD 39 334 VDD P12LL L=6E-08 W=8E-07 $X=4720 $Y=20545 $D=1
M467 70 9 VDD VDD P12LL L=6E-08 W=6E-07 $X=4730 $Y=8205 $D=1
M468 71 10 VDD VDD P12LL L=6E-08 W=6E-07 $X=4730 $Y=24890 $D=1
M469 VDD 65 102 VDD P12LL L=6E-08 W=8E-07 $X=4840 $Y=17355 $D=1
M470 VDD 61 LBLX[4] VDD P12LL L=6E-08 W=1E-06 $X=5005 $Y=1635 $D=1
M471 VDD 62 UBLX[4] VDD P12LL L=6E-08 W=1E-06 $X=5005 $Y=31060 $D=1
M472 VDD 72 70 VDD P12LL L=6E-08 W=6E-07 $X=5010 $Y=8205 $D=1
M473 335 35 VDD VDD P12LL L=6E-08 W=8E-07 $X=5010 $Y=13360 $D=1
M474 336 39 VDD VDD P12LL L=6E-08 W=8E-07 $X=5010 $Y=20545 $D=1
M475 VDD 72 71 VDD P12LL L=6E-08 W=6E-07 $X=5010 $Y=24890 $D=1
M476 26 9 335 VDD P12LL L=6E-08 W=8E-07 $X=5300 $Y=13360 $D=1
M477 27 10 336 VDD P12LL L=6E-08 W=8E-07 $X=5300 $Y=20545 $D=1
M478 80 72 VDD VDD P12LL L=6E-08 W=6E-07 $X=5430 $Y=8205 $D=1
M479 81 72 VDD VDD P12LL L=6E-08 W=6E-07 $X=5430 $Y=24890 $D=1
M480 LBLX[5] 82 VDD VDD P12LL L=6E-08 W=1E-06 $X=5435 $Y=1635 $D=1
M481 UBLX[5] 83 VDD VDD P12LL L=6E-08 W=1E-06 $X=5435 $Y=31060 $D=1
M482 72 YX[2] VDD VDD P12LL L=6E-08 W=4E-07 $X=5580 $Y=22045 $D=1
M483 VDD YX[2] 72 VDD P12LL L=6E-08 W=4E-07 $X=5580 $Y=22315 $D=1
M484 72 YX[2] VDD VDD P12LL L=6E-08 W=4E-07 $X=5580 $Y=22585 $D=1
M485 VDD 26 80 VDD P12LL L=6E-08 W=6E-07 $X=5710 $Y=8205 $D=1
M486 VDD 27 81 VDD P12LL L=6E-08 W=6E-07 $X=5710 $Y=24890 $D=1
M487 LBL[5] 82 LBLX[5] VDD P12LL L=6E-08 W=1E-06 $X=5745 $Y=1635 $D=1
M488 UBL[5] 83 UBLX[5] VDD P12LL L=6E-08 W=1E-06 $X=5745 $Y=31060 $D=1
M489 LBLX[5] 80 122 VDD P12LL L=6E-08 W=6E-07 $X=5945 $Y=5965 $D=1
M490 LBL[5] 80 110 VDD P12LL L=6E-08 W=6E-07 $X=5945 $Y=6885 $D=1
M491 UBL[5] 81 110 VDD P12LL L=6E-08 W=6E-07 $X=5945 $Y=26210 $D=1
M492 UBLX[5] 81 122 VDD P12LL L=6E-08 W=6E-07 $X=5945 $Y=27130 $D=1
M493 82 80 VDD VDD P12LL L=6E-08 W=6E-07 $X=5990 $Y=8205 $D=1
M494 83 81 VDD VDD P12LL L=6E-08 W=6E-07 $X=5990 $Y=24890 $D=1
M495 VDD 82 LBL[5] VDD P12LL L=6E-08 W=1E-06 $X=6055 $Y=1635 $D=1
M496 VDD 83 UBL[5] VDD P12LL L=6E-08 W=1E-06 $X=6055 $Y=31060 $D=1
M497 LBL[7] 84 VDD VDD P12LL L=6E-08 W=1E-06 $X=6485 $Y=1635 $D=1
M498 UBL[7] 85 VDD VDD P12LL L=6E-08 W=1E-06 $X=6485 $Y=31060 $D=1
M499 VDD 92 84 VDD P12LL L=6E-08 W=6E-07 $X=6550 $Y=8205 $D=1
M500 VDD 93 85 VDD P12LL L=6E-08 W=6E-07 $X=6550 $Y=24890 $D=1
M501 VDD 111 DOUT VDD P12LL L=6E-08 W=1E-06 $X=6585 $Y=13265 $D=1
M502 122 92 LBLX[7] VDD P12LL L=6E-08 W=6E-07 $X=6595 $Y=5965 $D=1
M503 110 92 LBL[7] VDD P12LL L=6E-08 W=6E-07 $X=6595 $Y=6885 $D=1
M504 110 93 UBL[7] VDD P12LL L=6E-08 W=6E-07 $X=6595 $Y=26210 $D=1
M505 122 93 UBLX[7] VDD P12LL L=6E-08 W=6E-07 $X=6595 $Y=27130 $D=1
M506 94 YX[3] VDD VDD P12LL L=6E-08 W=4E-07 $X=6620 $Y=22045 $D=1
M507 VDD YX[3] 94 VDD P12LL L=6E-08 W=4E-07 $X=6620 $Y=22315 $D=1
M508 94 YX[3] VDD VDD P12LL L=6E-08 W=4E-07 $X=6620 $Y=22585 $D=1
M509 LBLX[7] 84 LBL[7] VDD P12LL L=6E-08 W=1E-06 $X=6795 $Y=1635 $D=1
M510 UBLX[7] 85 UBL[7] VDD P12LL L=6E-08 W=1E-06 $X=6795 $Y=31060 $D=1
M511 92 26 VDD VDD P12LL L=6E-08 W=6E-07 $X=6830 $Y=8205 $D=1
M512 93 27 VDD VDD P12LL L=6E-08 W=6E-07 $X=6830 $Y=24890 $D=1
M513 DOUT 111 VDD VDD P12LL L=6E-08 W=1E-06 $X=6875 $Y=13265 $D=1
M514 VDD 84 LBLX[7] VDD P12LL L=6E-08 W=1E-06 $X=7105 $Y=1635 $D=1
M515 VDD 85 UBLX[7] VDD P12LL L=6E-08 W=1E-06 $X=7105 $Y=31060 $D=1
M516 VDD 94 92 VDD P12LL L=6E-08 W=6E-07 $X=7110 $Y=8205 $D=1
M517 VDD 94 93 VDD P12LL L=6E-08 W=6E-07 $X=7110 $Y=24890 $D=1
M518 VDD 111 DOUT VDD P12LL L=6E-08 W=1E-06 $X=7165 $Y=13265 $D=1
M519 105 94 VDD VDD P12LL L=6E-08 W=6E-07 $X=7530 $Y=8205 $D=1
M520 106 94 VDD VDD P12LL L=6E-08 W=6E-07 $X=7530 $Y=24890 $D=1
M521 LBLX[6] 107 VDD VDD P12LL L=6E-08 W=1E-06 $X=7535 $Y=1635 $D=1
M522 UBLX[6] 108 VDD VDD P12LL L=6E-08 W=1E-06 $X=7535 $Y=31060 $D=1
M523 103 109 110 VDD P12LL L=6E-08 W=7E-07 $X=7770 $Y=19600 $D=1
M524 103 116 VDD VDD P12LL L=1E-07 W=4E-07 $X=7795 $Y=18660 $D=1
M525 VDD 9 105 VDD P12LL L=6E-08 W=6E-07 $X=7810 $Y=8205 $D=1
M526 VDD 10 106 VDD P12LL L=6E-08 W=6E-07 $X=7810 $Y=24890 $D=1
M527 LBL[6] 107 LBLX[6] VDD P12LL L=6E-08 W=1E-06 $X=7845 $Y=1635 $D=1
M528 UBL[6] 108 UBLX[6] VDD P12LL L=6E-08 W=1E-06 $X=7845 $Y=31060 $D=1
M529 111 103 VDD VDD P12LL L=6E-08 W=1E-06 $X=7930 $Y=13160 $D=1
M530 LBLX[6] 105 122 VDD P12LL L=6E-08 W=6E-07 $X=8045 $Y=5965 $D=1
M531 LBL[6] 105 110 VDD P12LL L=6E-08 W=6E-07 $X=8045 $Y=6885 $D=1
M532 UBL[6] 106 110 VDD P12LL L=6E-08 W=6E-07 $X=8045 $Y=26210 $D=1
M533 UBLX[6] 106 122 VDD P12LL L=6E-08 W=6E-07 $X=8045 $Y=27130 $D=1
M534 110 109 103 VDD P12LL L=6E-08 W=7E-07 $X=8060 $Y=19600 $D=1
M535 110 102 VDD VDD P12LL L=6E-08 W=1E-06 $X=8080 $Y=20670 $D=1
M536 107 105 VDD VDD P12LL L=6E-08 W=6E-07 $X=8090 $Y=8205 $D=1
M537 108 106 VDD VDD P12LL L=6E-08 W=6E-07 $X=8090 $Y=24890 $D=1
M538 VDD 107 LBL[6] VDD P12LL L=6E-08 W=1E-06 $X=8155 $Y=1635 $D=1
M539 VDD 108 UBL[6] VDD P12LL L=6E-08 W=1E-06 $X=8155 $Y=31060 $D=1
M540 VDD 116 103 VDD P12LL L=1E-07 W=4E-07 $X=8165 $Y=18660 $D=1
M541 VDD 121 111 VDD P12LL L=6E-08 W=1E-06 $X=8220 $Y=13160 $D=1
M542 122 102 110 VDD P12LL L=6E-08 W=1E-06 $X=8370 $Y=20670 $D=1
M543 121 111 VDD VDD P12LL L=6E-08 W=1E-06 $X=8510 $Y=13160 $D=1
M544 116 103 VDD VDD P12LL L=1E-07 W=4E-07 $X=8535 $Y=18660 $D=1
M545 LBL[8] 112 VDD VDD P12LL L=6E-08 W=1E-06 $X=8585 $Y=1635 $D=1
M546 UBL[8] 113 VDD VDD P12LL L=6E-08 W=1E-06 $X=8585 $Y=31060 $D=1
M547 VDD 124 112 VDD P12LL L=6E-08 W=6E-07 $X=8650 $Y=8205 $D=1
M548 VDD 125 113 VDD P12LL L=6E-08 W=6E-07 $X=8650 $Y=24890 $D=1
M549 VDD 102 122 VDD P12LL L=6E-08 W=1E-06 $X=8660 $Y=20670 $D=1
M550 116 109 122 VDD P12LL L=6E-08 W=7E-07 $X=8680 $Y=19600 $D=1
M551 122 124 LBLX[8] VDD P12LL L=6E-08 W=6E-07 $X=8695 $Y=5965 $D=1
M552 110 124 LBL[8] VDD P12LL L=6E-08 W=6E-07 $X=8695 $Y=6885 $D=1
M553 110 125 UBL[8] VDD P12LL L=6E-08 W=6E-07 $X=8695 $Y=26210 $D=1
M554 122 125 UBLX[8] VDD P12LL L=6E-08 W=6E-07 $X=8695 $Y=27130 $D=1
M555 VDD 116 121 VDD P12LL L=6E-08 W=1E-06 $X=8800 $Y=13160 $D=1
M556 LBLX[8] 112 LBL[8] VDD P12LL L=6E-08 W=1E-06 $X=8895 $Y=1635 $D=1
M557 UBLX[8] 113 UBL[8] VDD P12LL L=6E-08 W=1E-06 $X=8895 $Y=31060 $D=1
M558 VDD 103 116 VDD P12LL L=1E-07 W=4E-07 $X=8905 $Y=18660 $D=1
M559 124 9 VDD VDD P12LL L=6E-08 W=6E-07 $X=8930 $Y=8205 $D=1
M560 125 10 VDD VDD P12LL L=6E-08 W=6E-07 $X=8930 $Y=24890 $D=1
M561 122 109 116 VDD P12LL L=6E-08 W=7E-07 $X=8970 $Y=19600 $D=1
M562 VDD 112 LBLX[8] VDD P12LL L=6E-08 W=1E-06 $X=9205 $Y=1635 $D=1
M563 VDD 113 UBLX[8] VDD P12LL L=6E-08 W=1E-06 $X=9205 $Y=31060 $D=1
M564 VDD 126 124 VDD P12LL L=6E-08 W=6E-07 $X=9210 $Y=8205 $D=1
M565 VDD 126 125 VDD P12LL L=6E-08 W=6E-07 $X=9210 $Y=24890 $D=1
M566 134 126 VDD VDD P12LL L=6E-08 W=6E-07 $X=9630 $Y=8205 $D=1
M567 135 126 VDD VDD P12LL L=6E-08 W=6E-07 $X=9630 $Y=24890 $D=1
M568 LBLX[9] 137 VDD VDD P12LL L=6E-08 W=1E-06 $X=9635 $Y=1635 $D=1
M569 UBLX[9] 138 VDD VDD P12LL L=6E-08 W=1E-06 $X=9635 $Y=31060 $D=1
M570 VDD YX[4] 126 VDD P12LL L=6E-08 W=4E-07 $X=9780 $Y=11050 $D=1
M571 126 YX[4] VDD VDD P12LL L=6E-08 W=4E-07 $X=9780 $Y=11320 $D=1
M572 VDD YX[4] 126 VDD P12LL L=6E-08 W=4E-07 $X=9780 $Y=11590 $D=1
M573 VDD 26 134 VDD P12LL L=6E-08 W=6E-07 $X=9910 $Y=8205 $D=1
M574 VDD 27 135 VDD P12LL L=6E-08 W=6E-07 $X=9910 $Y=24890 $D=1
M575 LBL[9] 137 LBLX[9] VDD P12LL L=6E-08 W=1E-06 $X=9945 $Y=1635 $D=1
M576 UBL[9] 138 UBLX[9] VDD P12LL L=6E-08 W=1E-06 $X=9945 $Y=31060 $D=1
M577 LBLX[9] 134 122 VDD P12LL L=6E-08 W=6E-07 $X=10145 $Y=5965 $D=1
M578 LBL[9] 134 110 VDD P12LL L=6E-08 W=6E-07 $X=10145 $Y=6885 $D=1
M579 UBL[9] 135 110 VDD P12LL L=6E-08 W=6E-07 $X=10145 $Y=26210 $D=1
M580 UBLX[9] 135 122 VDD P12LL L=6E-08 W=6E-07 $X=10145 $Y=27130 $D=1
M581 137 134 VDD VDD P12LL L=6E-08 W=6E-07 $X=10190 $Y=8205 $D=1
M582 138 135 VDD VDD P12LL L=6E-08 W=6E-07 $X=10190 $Y=24890 $D=1
M583 VDD DATA 140 VDD P12LL L=6E-08 W=4E-07 $X=10195 $Y=13885 $D=1
M584 VDD 137 LBL[9] VDD P12LL L=6E-08 W=1E-06 $X=10255 $Y=1635 $D=1
M585 VDD 138 UBL[9] VDD P12LL L=6E-08 W=1E-06 $X=10255 $Y=31060 $D=1
M586 150 140 VDD VDD P12LL L=3E-07 W=4E-07 $X=10545 $Y=13885 $D=1
M587 VDD 147 139 VDD P12LL L=6E-08 W=1E-06 $X=10590 $Y=20595 $D=1
M588 LBL[11] 141 VDD VDD P12LL L=6E-08 W=1E-06 $X=10685 $Y=1635 $D=1
M589 UBL[11] 142 VDD VDD P12LL L=6E-08 W=1E-06 $X=10685 $Y=31060 $D=1
M590 VDD 151 141 VDD P12LL L=6E-08 W=6E-07 $X=10750 $Y=8205 $D=1
M591 VDD 152 142 VDD P12LL L=6E-08 W=6E-07 $X=10750 $Y=24890 $D=1
M592 122 151 LBLX[11] VDD P12LL L=6E-08 W=6E-07 $X=10795 $Y=5965 $D=1
M593 110 151 LBL[11] VDD P12LL L=6E-08 W=6E-07 $X=10795 $Y=6885 $D=1
M594 110 152 UBL[11] VDD P12LL L=6E-08 W=6E-07 $X=10795 $Y=26210 $D=1
M595 122 152 UBLX[11] VDD P12LL L=6E-08 W=6E-07 $X=10795 $Y=27130 $D=1
M596 VDD YX[5] 153 VDD P12LL L=6E-08 W=4E-07 $X=10820 $Y=11050 $D=1
M597 153 YX[5] VDD VDD P12LL L=6E-08 W=4E-07 $X=10820 $Y=11320 $D=1
M598 VDD YX[5] 153 VDD P12LL L=6E-08 W=4E-07 $X=10820 $Y=11590 $D=1
M599 147 SACK1 VDD VDD P12LL L=6E-08 W=4E-07 $X=10890 $Y=20595 $D=1
M600 LBLX[11] 141 LBL[11] VDD P12LL L=6E-08 W=1E-06 $X=10995 $Y=1635 $D=1
M601 UBLX[11] 142 UBL[11] VDD P12LL L=6E-08 W=1E-06 $X=10995 $Y=31060 $D=1
M602 VDD VDD DATA VDD P12LL L=6E-08 W=2E-07 $X=11015 $Y=13170 $D=1
M603 151 26 VDD VDD P12LL L=6E-08 W=6E-07 $X=11030 $Y=8205 $D=1
M604 152 27 VDD VDD P12LL L=6E-08 W=6E-07 $X=11030 $Y=24890 $D=1
M605 VDD 141 LBLX[11] VDD P12LL L=6E-08 W=1E-06 $X=11305 $Y=1635 $D=1
M606 VDD 142 UBLX[11] VDD P12LL L=6E-08 W=1E-06 $X=11305 $Y=31060 $D=1
M607 VDD 153 151 VDD P12LL L=6E-08 W=6E-07 $X=11310 $Y=8205 $D=1
M608 VDD 153 152 VDD P12LL L=6E-08 W=6E-07 $X=11310 $Y=24890 $D=1
M609 VDD 202 185 VDD P12LL L=6E-08 W=4E-07 $X=11405 $Y=17435 $D=1
M610 VDD 150 159 VDD P12LL L=2E-07 W=4E-07 $X=11505 $Y=13885 $D=1
M611 VDD 165 109 VDD P12LL L=6E-08 W=1E-06 $X=11515 $Y=20595 $D=1
M612 163 153 VDD VDD P12LL L=6E-08 W=6E-07 $X=11730 $Y=8205 $D=1
M613 164 153 VDD VDD P12LL L=6E-08 W=6E-07 $X=11730 $Y=24890 $D=1
M614 LBLX[10] 166 VDD VDD P12LL L=6E-08 W=1E-06 $X=11735 $Y=1635 $D=1
M615 UBLX[10] 167 VDD VDD P12LL L=6E-08 W=1E-06 $X=11735 $Y=31060 $D=1
M616 165 SACK1 VDD VDD P12LL L=6E-08 W=4E-07 $X=11815 $Y=20595 $D=1
M617 168 159 VDD VDD P12LL L=6E-08 W=7E-07 $X=11995 $Y=13585 $D=1
M618 VDD 9 163 VDD P12LL L=6E-08 W=6E-07 $X=12010 $Y=8205 $D=1
M619 VDD 10 164 VDD P12LL L=6E-08 W=6E-07 $X=12010 $Y=24890 $D=1
M620 LBL[10] 166 LBLX[10] VDD P12LL L=6E-08 W=1E-06 $X=12045 $Y=1635 $D=1
M621 UBL[10] 167 UBLX[10] VDD P12LL L=6E-08 W=1E-06 $X=12045 $Y=31060 $D=1
M622 VDD SACK4 165 VDD P12LL L=6E-08 W=4E-07 $X=12105 $Y=20595 $D=1
M623 LBLX[10] 163 122 VDD P12LL L=6E-08 W=6E-07 $X=12245 $Y=5965 $D=1
M624 LBL[10] 163 110 VDD P12LL L=6E-08 W=6E-07 $X=12245 $Y=6885 $D=1
M625 UBL[10] 164 110 VDD P12LL L=6E-08 W=6E-07 $X=12245 $Y=26210 $D=1
M626 UBLX[10] 164 122 VDD P12LL L=6E-08 W=6E-07 $X=12245 $Y=27130 $D=1
M627 166 163 VDD VDD P12LL L=6E-08 W=6E-07 $X=12290 $Y=8205 $D=1
M628 167 164 VDD VDD P12LL L=6E-08 W=6E-07 $X=12290 $Y=24890 $D=1
M629 VDD 166 LBL[10] VDD P12LL L=6E-08 W=1E-06 $X=12355 $Y=1635 $D=1
M630 VDD 167 UBL[10] VDD P12LL L=6E-08 W=1E-06 $X=12355 $Y=31060 $D=1
M631 VDD 202 172 VDD P12LL L=3E-07 W=1.2E-07 $X=12455 $Y=17335 $D=1
M632 169 193 VDD VDD P12LL L=6E-08 W=1E-06 $X=12460 $Y=20595 $D=1
M633 172 CLK 168 VDD P12LL L=6E-08 W=7E-07 $X=12675 $Y=13695 $D=1
M634 VDD 193 169 VDD P12LL L=6E-08 W=1E-06 $X=12750 $Y=20595 $D=1
M635 LBL[12] 173 VDD VDD P12LL L=6E-08 W=1E-06 $X=12785 $Y=1635 $D=1
M636 UBL[12] 174 VDD VDD P12LL L=6E-08 W=1E-06 $X=12785 $Y=31060 $D=1
M637 VDD 181 173 VDD P12LL L=6E-08 W=6E-07 $X=12850 $Y=8205 $D=1
M638 VDD 182 174 VDD P12LL L=6E-08 W=6E-07 $X=12850 $Y=24890 $D=1
M639 122 181 LBLX[12] VDD P12LL L=6E-08 W=6E-07 $X=12895 $Y=5965 $D=1
M640 110 181 LBL[12] VDD P12LL L=6E-08 W=6E-07 $X=12895 $Y=6885 $D=1
M641 110 182 UBL[12] VDD P12LL L=6E-08 W=6E-07 $X=12895 $Y=26210 $D=1
M642 122 182 UBLX[12] VDD P12LL L=6E-08 W=6E-07 $X=12895 $Y=27130 $D=1
M643 169 193 VDD VDD P12LL L=6E-08 W=1E-06 $X=13040 $Y=20595 $D=1
M644 202 172 VDD VDD P12LL L=6E-08 W=8E-07 $X=13090 $Y=17335 $D=1
M645 LBLX[12] 173 LBL[12] VDD P12LL L=6E-08 W=1E-06 $X=13095 $Y=1635 $D=1
M646 UBLX[12] 174 UBL[12] VDD P12LL L=6E-08 W=1E-06 $X=13095 $Y=31060 $D=1
M647 181 9 VDD VDD P12LL L=6E-08 W=6E-07 $X=13130 $Y=8205 $D=1
M648 182 10 VDD VDD P12LL L=6E-08 W=6E-07 $X=13130 $Y=24890 $D=1
M649 188 CLK 200 VDD P12LL L=6E-08 W=7E-07 $X=13295 $Y=13695 $D=1
M650 VDD 193 169 VDD P12LL L=6E-08 W=1E-06 $X=13330 $Y=20595 $D=1
M651 VDD 173 LBLX[12] VDD P12LL L=6E-08 W=1E-06 $X=13405 $Y=1635 $D=1
M652 VDD 174 UBLX[12] VDD P12LL L=6E-08 W=1E-06 $X=13405 $Y=31060 $D=1
M653 VDD 183 181 VDD P12LL L=6E-08 W=6E-07 $X=13410 $Y=8205 $D=1
M654 VDD 183 182 VDD P12LL L=6E-08 W=6E-07 $X=13410 $Y=24890 $D=1
M655 193 185 VDD VDD P12LL L=6E-08 W=8E-07 $X=13620 $Y=20595 $D=1
M656 VDD 200 212 VDD P12LL L=6E-08 W=4E-07 $X=13750 $Y=17335 $D=1
M657 194 183 VDD VDD P12LL L=6E-08 W=6E-07 $X=13830 $Y=8205 $D=1
M658 195 183 VDD VDD P12LL L=6E-08 W=6E-07 $X=13830 $Y=24890 $D=1
M659 LBLX[13] 196 VDD VDD P12LL L=6E-08 W=1E-06 $X=13835 $Y=1635 $D=1
M660 UBLX[13] 197 VDD VDD P12LL L=6E-08 W=1E-06 $X=13835 $Y=31060 $D=1
M661 VDD 227 193 VDD P12LL L=6E-08 W=8E-07 $X=13925 $Y=20595 $D=1
M662 VDD 198 188 VDD P12LL L=6E-08 W=7E-07 $X=13955 $Y=13585 $D=1
M663 VDD YX[6] 183 VDD P12LL L=6E-08 W=4E-07 $X=13980 $Y=11050 $D=1
M664 183 YX[6] VDD VDD P12LL L=6E-08 W=4E-07 $X=13980 $Y=11320 $D=1
M665 VDD YX[6] 183 VDD P12LL L=6E-08 W=4E-07 $X=13980 $Y=11590 $D=1
M666 VDD 26 194 VDD P12LL L=6E-08 W=6E-07 $X=14110 $Y=8205 $D=1
M667 VDD 27 195 VDD P12LL L=6E-08 W=6E-07 $X=14110 $Y=24890 $D=1
M668 LBL[13] 196 LBLX[13] VDD P12LL L=6E-08 W=1E-06 $X=14145 $Y=1635 $D=1
M669 200 212 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=14145 $Y=17335 $D=1
M670 UBL[13] 197 UBLX[13] VDD P12LL L=6E-08 W=1E-06 $X=14145 $Y=31060 $D=1
M671 198 207 VDD VDD P12LL L=2E-07 W=4E-07 $X=14305 $Y=13885 $D=1
M672 LBLX[13] 194 122 VDD P12LL L=6E-08 W=6E-07 $X=14345 $Y=5965 $D=1
M673 LBL[13] 194 110 VDD P12LL L=6E-08 W=6E-07 $X=14345 $Y=6885 $D=1
M674 UBL[13] 195 110 VDD P12LL L=6E-08 W=6E-07 $X=14345 $Y=26210 $D=1
M675 UBLX[13] 195 122 VDD P12LL L=6E-08 W=6E-07 $X=14345 $Y=27130 $D=1
M676 196 194 VDD VDD P12LL L=6E-08 W=6E-07 $X=14390 $Y=8205 $D=1
M677 197 195 VDD VDD P12LL L=6E-08 W=6E-07 $X=14390 $Y=24890 $D=1
M678 VDD 196 LBL[13] VDD P12LL L=6E-08 W=1E-06 $X=14455 $Y=1635 $D=1
M679 VDD 197 UBL[13] VDD P12LL L=6E-08 W=1E-06 $X=14455 $Y=31060 $D=1
M680 201 227 VDD VDD P12LL L=6E-08 W=8E-07 $X=14605 $Y=20595 $D=1
M681 LBL[15] 203 VDD VDD P12LL L=6E-08 W=1E-06 $X=14885 $Y=1635 $D=1
M682 UBL[15] 204 VDD VDD P12LL L=6E-08 W=1E-06 $X=14885 $Y=31060 $D=1
M683 VDD 202 201 VDD P12LL L=6E-08 W=8E-07 $X=14910 $Y=20595 $D=1
M684 VDD 213 203 VDD P12LL L=6E-08 W=6E-07 $X=14950 $Y=8205 $D=1
M685 VDD 215 204 VDD P12LL L=6E-08 W=6E-07 $X=14950 $Y=24890 $D=1
M686 122 213 LBLX[15] VDD P12LL L=6E-08 W=6E-07 $X=14995 $Y=5965 $D=1
M687 110 213 LBL[15] VDD P12LL L=6E-08 W=6E-07 $X=14995 $Y=6885 $D=1
M688 110 215 UBL[15] VDD P12LL L=6E-08 W=6E-07 $X=14995 $Y=26210 $D=1
M689 122 215 UBLX[15] VDD P12LL L=6E-08 W=6E-07 $X=14995 $Y=27130 $D=1
M690 VDD YX[7] 214 VDD P12LL L=6E-08 W=4E-07 $X=15020 $Y=11050 $D=1
M691 214 YX[7] VDD VDD P12LL L=6E-08 W=4E-07 $X=15020 $Y=11320 $D=1
M692 VDD YX[7] 214 VDD P12LL L=6E-08 W=4E-07 $X=15020 $Y=11590 $D=1
M693 VDD 217 207 VDD P12LL L=3E-07 W=4E-07 $X=15165 $Y=13885 $D=1
M694 LBLX[15] 203 LBL[15] VDD P12LL L=6E-08 W=1E-06 $X=15195 $Y=1635 $D=1
M695 UBLX[15] 204 UBL[15] VDD P12LL L=6E-08 W=1E-06 $X=15195 $Y=31060 $D=1
M696 199 201 VDD VDD P12LL L=6E-08 W=1E-06 $X=15200 $Y=20595 $D=1
M697 213 26 VDD VDD P12LL L=6E-08 W=6E-07 $X=15230 $Y=8205 $D=1
M698 215 27 VDD VDD P12LL L=6E-08 W=6E-07 $X=15230 $Y=24890 $D=1
M699 220 212 VDD VDD P12LL L=6E-08 W=4E-07 $X=15460 $Y=17295 $D=1
M700 VDD 201 199 VDD P12LL L=6E-08 W=1E-06 $X=15490 $Y=20595 $D=1
M701 VDD 203 LBLX[15] VDD P12LL L=6E-08 W=1E-06 $X=15505 $Y=1635 $D=1
M702 VDD 204 UBLX[15] VDD P12LL L=6E-08 W=1E-06 $X=15505 $Y=31060 $D=1
M703 VDD 214 213 VDD P12LL L=6E-08 W=6E-07 $X=15510 $Y=8205 $D=1
M704 VDD 214 215 VDD P12LL L=6E-08 W=6E-07 $X=15510 $Y=24890 $D=1
M705 217 226 VDD VDD P12LL L=6E-08 W=4E-07 $X=15755 $Y=13885 $D=1
M706 VDD WE 220 VDD P12LL L=6E-08 W=4E-07 $X=15765 $Y=17295 $D=1
M707 199 201 VDD VDD P12LL L=6E-08 W=1E-06 $X=15780 $Y=20595 $D=1
M708 228 214 VDD VDD P12LL L=6E-08 W=6E-07 $X=15930 $Y=8205 $D=1
M709 229 214 VDD VDD P12LL L=6E-08 W=6E-07 $X=15930 $Y=24890 $D=1
M710 LBLX[14] 231 VDD VDD P12LL L=6E-08 W=1E-06 $X=15935 $Y=1635 $D=1
M711 UBLX[14] 232 VDD VDD P12LL L=6E-08 W=1E-06 $X=15935 $Y=31060 $D=1
M712 227 220 VDD VDD P12LL L=6E-08 W=1E-06 $X=16055 $Y=17295 $D=1
M713 VDD 201 199 VDD P12LL L=6E-08 W=1E-06 $X=16070 $Y=20595 $D=1
M714 230 230 VDD VDD P12LL L=6E-08 W=4E-07 $X=16190 $Y=13085 $D=1
M715 VDD 9 228 VDD P12LL L=6E-08 W=6E-07 $X=16210 $Y=8205 $D=1
M716 VDD 10 229 VDD P12LL L=6E-08 W=6E-07 $X=16210 $Y=24890 $D=1
M717 LBL[14] 231 LBLX[14] VDD P12LL L=6E-08 W=1E-06 $X=16245 $Y=1635 $D=1
M718 UBL[14] 232 UBLX[14] VDD P12LL L=6E-08 W=1E-06 $X=16245 $Y=31060 $D=1
M719 LBLX[14] 228 122 VDD P12LL L=6E-08 W=6E-07 $X=16445 $Y=5965 $D=1
M720 LBL[14] 228 110 VDD P12LL L=6E-08 W=6E-07 $X=16445 $Y=6885 $D=1
M721 UBL[14] 229 110 VDD P12LL L=6E-08 W=6E-07 $X=16445 $Y=26210 $D=1
M722 UBLX[14] 229 122 VDD P12LL L=6E-08 W=6E-07 $X=16445 $Y=27130 $D=1
M723 231 228 VDD VDD P12LL L=6E-08 W=6E-07 $X=16490 $Y=8205 $D=1
M724 232 229 VDD VDD P12LL L=6E-08 W=6E-07 $X=16490 $Y=24890 $D=1
M725 VDD 231 LBL[14] VDD P12LL L=6E-08 W=1E-06 $X=16555 $Y=1635 $D=1
M726 VDD 232 UBL[14] VDD P12LL L=6E-08 W=1E-06 $X=16555 $Y=31060 $D=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_Y16_X512_D1
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_Y16_X512_D1 D[0] DCTRCLK DCTRCLKX Q[0] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX
XI0 LBL[15] LBL[14] LBLX[15] LBLX[14] STWL RWLL[0] RWLL[1] VDD VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN
XI1 LBL[13] LBL[12] LBLX[13] LBLX[12] STWL RWLL[0] RWLL[1] VDD VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN
XI2 LBL[11] LBL[10] LBLX[11] LBLX[10] STWL RWLL[0] RWLL[1] VDD VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN
XI3 LBL[9] LBL[8] LBLX[9] LBLX[8] STWL RWLL[0] RWLL[1] VDD VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN
XI4 LBL[7] LBL[6] LBLX[7] LBLX[6] STWL RWLL[0] RWLL[1] VDD VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN
XI5 LBL[5] LBL[4] LBLX[5] LBLX[4] STWL RWLL[0] RWLL[1] VDD VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN
XI6 LBL[3] LBL[2] LBLX[3] LBLX[2] STWL RWLL[0] RWLL[1] VDD VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN
XI7 LBL[1] LBL[0] LBLX[1] LBLX[0] STWL RWLL[0] RWLL[1] VDD VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN
XI8 UBL[15] UBL[14] UBLX[15] UBLX[14] RWLU[0] RWLU[1] VDD VSS WL[511] WL[510]
+WL[509] WL[508] WL[507] WL[506] WL[505] WL[504] WL[503] WL[502] WL[501] WL[500]
+WL[499] WL[498] WL[497] WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] WL[490]
+WL[489] WL[488] WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480]
+WL[479] WL[478] WL[477] WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] WL[470]
+WL[469] WL[468] WL[467] WL[466] WL[465] WL[464] WL[463] WL[462] WL[461] WL[460]
+WL[459] WL[458] WL[457] WL[456] WL[455] WL[454] WL[453] WL[452] WL[451] WL[450]
+WL[449] WL[448] WL[447] WL[446] WL[445] WL[444] WL[443] WL[442] WL[441] WL[440]
+WL[439] WL[438] WL[437] WL[436] WL[435] WL[434] WL[433] WL[432] WL[431] WL[430]
+WL[429] WL[428] WL[427] WL[426] WL[425] WL[424] WL[423] WL[422] WL[421] WL[420]
+WL[419] WL[418] WL[417] WL[416] WL[415] WL[414] WL[413] WL[412] WL[411] WL[410]
+WL[409] WL[408] WL[407] WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] WL[400]
+WL[399] WL[398] WL[397] WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390]
+WL[389] WL[388] WL[387] WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] WL[380]
+WL[379] WL[378] WL[377] WL[376] WL[375] WL[374] WL[373] WL[372] WL[371] WL[370]
+WL[369] WL[368] WL[367] WL[366] WL[365] WL[364] WL[363] WL[362] WL[361] WL[360]
+WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] WL[353] WL[352] WL[351] WL[350]
+WL[349] WL[348] WL[347] WL[346] WL[345] WL[344] WL[343] WL[342] WL[341] WL[340]
+WL[339] WL[338] WL[337] WL[336] WL[335] WL[334] WL[333] WL[332] WL[331] WL[330]
+WL[329] WL[328] WL[327] WL[326] WL[325] WL[324] WL[323] WL[322] WL[321] WL[320]
+WL[319] WL[318] WL[317] WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] WL[310]
+WL[309] WL[308] WL[307] WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300]
+WL[299] WL[298] WL[297] WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] WL[290]
+WL[289] WL[288] WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] WL[281] WL[280]
+WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273] WL[272] WL[271] WL[270]
+WL[269] WL[268] WL[267] WL[266] WL[265] WL[264] WL[263] WL[262] WL[261] WL[260]
+WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_UP
XI9 UBL[13] UBL[12] UBLX[13] UBLX[12] RWLU[0] RWLU[1] VDD VSS WL[511] WL[510]
+WL[509] WL[508] WL[507] WL[506] WL[505] WL[504] WL[503] WL[502] WL[501] WL[500]
+WL[499] WL[498] WL[497] WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] WL[490]
+WL[489] WL[488] WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480]
+WL[479] WL[478] WL[477] WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] WL[470]
+WL[469] WL[468] WL[467] WL[466] WL[465] WL[464] WL[463] WL[462] WL[461] WL[460]
+WL[459] WL[458] WL[457] WL[456] WL[455] WL[454] WL[453] WL[452] WL[451] WL[450]
+WL[449] WL[448] WL[447] WL[446] WL[445] WL[444] WL[443] WL[442] WL[441] WL[440]
+WL[439] WL[438] WL[437] WL[436] WL[435] WL[434] WL[433] WL[432] WL[431] WL[430]
+WL[429] WL[428] WL[427] WL[426] WL[425] WL[424] WL[423] WL[422] WL[421] WL[420]
+WL[419] WL[418] WL[417] WL[416] WL[415] WL[414] WL[413] WL[412] WL[411] WL[410]
+WL[409] WL[408] WL[407] WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] WL[400]
+WL[399] WL[398] WL[397] WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390]
+WL[389] WL[388] WL[387] WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] WL[380]
+WL[379] WL[378] WL[377] WL[376] WL[375] WL[374] WL[373] WL[372] WL[371] WL[370]
+WL[369] WL[368] WL[367] WL[366] WL[365] WL[364] WL[363] WL[362] WL[361] WL[360]
+WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] WL[353] WL[352] WL[351] WL[350]
+WL[349] WL[348] WL[347] WL[346] WL[345] WL[344] WL[343] WL[342] WL[341] WL[340]
+WL[339] WL[338] WL[337] WL[336] WL[335] WL[334] WL[333] WL[332] WL[331] WL[330]
+WL[329] WL[328] WL[327] WL[326] WL[325] WL[324] WL[323] WL[322] WL[321] WL[320]
+WL[319] WL[318] WL[317] WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] WL[310]
+WL[309] WL[308] WL[307] WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300]
+WL[299] WL[298] WL[297] WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] WL[290]
+WL[289] WL[288] WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] WL[281] WL[280]
+WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273] WL[272] WL[271] WL[270]
+WL[269] WL[268] WL[267] WL[266] WL[265] WL[264] WL[263] WL[262] WL[261] WL[260]
+WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_UP
XI10 UBL[11] UBL[10] UBLX[11] UBLX[10] RWLU[0] RWLU[1] VDD VSS WL[511] WL[510]
+WL[509] WL[508] WL[507] WL[506] WL[505] WL[504] WL[503] WL[502] WL[501] WL[500]
+WL[499] WL[498] WL[497] WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] WL[490]
+WL[489] WL[488] WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480]
+WL[479] WL[478] WL[477] WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] WL[470]
+WL[469] WL[468] WL[467] WL[466] WL[465] WL[464] WL[463] WL[462] WL[461] WL[460]
+WL[459] WL[458] WL[457] WL[456] WL[455] WL[454] WL[453] WL[452] WL[451] WL[450]
+WL[449] WL[448] WL[447] WL[446] WL[445] WL[444] WL[443] WL[442] WL[441] WL[440]
+WL[439] WL[438] WL[437] WL[436] WL[435] WL[434] WL[433] WL[432] WL[431] WL[430]
+WL[429] WL[428] WL[427] WL[426] WL[425] WL[424] WL[423] WL[422] WL[421] WL[420]
+WL[419] WL[418] WL[417] WL[416] WL[415] WL[414] WL[413] WL[412] WL[411] WL[410]
+WL[409] WL[408] WL[407] WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] WL[400]
+WL[399] WL[398] WL[397] WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390]
+WL[389] WL[388] WL[387] WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] WL[380]
+WL[379] WL[378] WL[377] WL[376] WL[375] WL[374] WL[373] WL[372] WL[371] WL[370]
+WL[369] WL[368] WL[367] WL[366] WL[365] WL[364] WL[363] WL[362] WL[361] WL[360]
+WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] WL[353] WL[352] WL[351] WL[350]
+WL[349] WL[348] WL[347] WL[346] WL[345] WL[344] WL[343] WL[342] WL[341] WL[340]
+WL[339] WL[338] WL[337] WL[336] WL[335] WL[334] WL[333] WL[332] WL[331] WL[330]
+WL[329] WL[328] WL[327] WL[326] WL[325] WL[324] WL[323] WL[322] WL[321] WL[320]
+WL[319] WL[318] WL[317] WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] WL[310]
+WL[309] WL[308] WL[307] WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300]
+WL[299] WL[298] WL[297] WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] WL[290]
+WL[289] WL[288] WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] WL[281] WL[280]
+WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273] WL[272] WL[271] WL[270]
+WL[269] WL[268] WL[267] WL[266] WL[265] WL[264] WL[263] WL[262] WL[261] WL[260]
+WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_UP
XI11 UBL[9] UBL[8] UBLX[9] UBLX[8] RWLU[0] RWLU[1] VDD VSS WL[511] WL[510]
+WL[509] WL[508] WL[507] WL[506] WL[505] WL[504] WL[503] WL[502] WL[501] WL[500]
+WL[499] WL[498] WL[497] WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] WL[490]
+WL[489] WL[488] WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480]
+WL[479] WL[478] WL[477] WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] WL[470]
+WL[469] WL[468] WL[467] WL[466] WL[465] WL[464] WL[463] WL[462] WL[461] WL[460]
+WL[459] WL[458] WL[457] WL[456] WL[455] WL[454] WL[453] WL[452] WL[451] WL[450]
+WL[449] WL[448] WL[447] WL[446] WL[445] WL[444] WL[443] WL[442] WL[441] WL[440]
+WL[439] WL[438] WL[437] WL[436] WL[435] WL[434] WL[433] WL[432] WL[431] WL[430]
+WL[429] WL[428] WL[427] WL[426] WL[425] WL[424] WL[423] WL[422] WL[421] WL[420]
+WL[419] WL[418] WL[417] WL[416] WL[415] WL[414] WL[413] WL[412] WL[411] WL[410]
+WL[409] WL[408] WL[407] WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] WL[400]
+WL[399] WL[398] WL[397] WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390]
+WL[389] WL[388] WL[387] WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] WL[380]
+WL[379] WL[378] WL[377] WL[376] WL[375] WL[374] WL[373] WL[372] WL[371] WL[370]
+WL[369] WL[368] WL[367] WL[366] WL[365] WL[364] WL[363] WL[362] WL[361] WL[360]
+WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] WL[353] WL[352] WL[351] WL[350]
+WL[349] WL[348] WL[347] WL[346] WL[345] WL[344] WL[343] WL[342] WL[341] WL[340]
+WL[339] WL[338] WL[337] WL[336] WL[335] WL[334] WL[333] WL[332] WL[331] WL[330]
+WL[329] WL[328] WL[327] WL[326] WL[325] WL[324] WL[323] WL[322] WL[321] WL[320]
+WL[319] WL[318] WL[317] WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] WL[310]
+WL[309] WL[308] WL[307] WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300]
+WL[299] WL[298] WL[297] WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] WL[290]
+WL[289] WL[288] WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] WL[281] WL[280]
+WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273] WL[272] WL[271] WL[270]
+WL[269] WL[268] WL[267] WL[266] WL[265] WL[264] WL[263] WL[262] WL[261] WL[260]
+WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_UP
XI12 UBL[7] UBL[6] UBLX[7] UBLX[6] RWLU[0] RWLU[1] VDD VSS WL[511] WL[510]
+WL[509] WL[508] WL[507] WL[506] WL[505] WL[504] WL[503] WL[502] WL[501] WL[500]
+WL[499] WL[498] WL[497] WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] WL[490]
+WL[489] WL[488] WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480]
+WL[479] WL[478] WL[477] WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] WL[470]
+WL[469] WL[468] WL[467] WL[466] WL[465] WL[464] WL[463] WL[462] WL[461] WL[460]
+WL[459] WL[458] WL[457] WL[456] WL[455] WL[454] WL[453] WL[452] WL[451] WL[450]
+WL[449] WL[448] WL[447] WL[446] WL[445] WL[444] WL[443] WL[442] WL[441] WL[440]
+WL[439] WL[438] WL[437] WL[436] WL[435] WL[434] WL[433] WL[432] WL[431] WL[430]
+WL[429] WL[428] WL[427] WL[426] WL[425] WL[424] WL[423] WL[422] WL[421] WL[420]
+WL[419] WL[418] WL[417] WL[416] WL[415] WL[414] WL[413] WL[412] WL[411] WL[410]
+WL[409] WL[408] WL[407] WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] WL[400]
+WL[399] WL[398] WL[397] WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390]
+WL[389] WL[388] WL[387] WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] WL[380]
+WL[379] WL[378] WL[377] WL[376] WL[375] WL[374] WL[373] WL[372] WL[371] WL[370]
+WL[369] WL[368] WL[367] WL[366] WL[365] WL[364] WL[363] WL[362] WL[361] WL[360]
+WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] WL[353] WL[352] WL[351] WL[350]
+WL[349] WL[348] WL[347] WL[346] WL[345] WL[344] WL[343] WL[342] WL[341] WL[340]
+WL[339] WL[338] WL[337] WL[336] WL[335] WL[334] WL[333] WL[332] WL[331] WL[330]
+WL[329] WL[328] WL[327] WL[326] WL[325] WL[324] WL[323] WL[322] WL[321] WL[320]
+WL[319] WL[318] WL[317] WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] WL[310]
+WL[309] WL[308] WL[307] WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300]
+WL[299] WL[298] WL[297] WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] WL[290]
+WL[289] WL[288] WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] WL[281] WL[280]
+WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273] WL[272] WL[271] WL[270]
+WL[269] WL[268] WL[267] WL[266] WL[265] WL[264] WL[263] WL[262] WL[261] WL[260]
+WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_UP
XI13 UBL[5] UBL[4] UBLX[5] UBLX[4] RWLU[0] RWLU[1] VDD VSS WL[511] WL[510]
+WL[509] WL[508] WL[507] WL[506] WL[505] WL[504] WL[503] WL[502] WL[501] WL[500]
+WL[499] WL[498] WL[497] WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] WL[490]
+WL[489] WL[488] WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480]
+WL[479] WL[478] WL[477] WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] WL[470]
+WL[469] WL[468] WL[467] WL[466] WL[465] WL[464] WL[463] WL[462] WL[461] WL[460]
+WL[459] WL[458] WL[457] WL[456] WL[455] WL[454] WL[453] WL[452] WL[451] WL[450]
+WL[449] WL[448] WL[447] WL[446] WL[445] WL[444] WL[443] WL[442] WL[441] WL[440]
+WL[439] WL[438] WL[437] WL[436] WL[435] WL[434] WL[433] WL[432] WL[431] WL[430]
+WL[429] WL[428] WL[427] WL[426] WL[425] WL[424] WL[423] WL[422] WL[421] WL[420]
+WL[419] WL[418] WL[417] WL[416] WL[415] WL[414] WL[413] WL[412] WL[411] WL[410]
+WL[409] WL[408] WL[407] WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] WL[400]
+WL[399] WL[398] WL[397] WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390]
+WL[389] WL[388] WL[387] WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] WL[380]
+WL[379] WL[378] WL[377] WL[376] WL[375] WL[374] WL[373] WL[372] WL[371] WL[370]
+WL[369] WL[368] WL[367] WL[366] WL[365] WL[364] WL[363] WL[362] WL[361] WL[360]
+WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] WL[353] WL[352] WL[351] WL[350]
+WL[349] WL[348] WL[347] WL[346] WL[345] WL[344] WL[343] WL[342] WL[341] WL[340]
+WL[339] WL[338] WL[337] WL[336] WL[335] WL[334] WL[333] WL[332] WL[331] WL[330]
+WL[329] WL[328] WL[327] WL[326] WL[325] WL[324] WL[323] WL[322] WL[321] WL[320]
+WL[319] WL[318] WL[317] WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] WL[310]
+WL[309] WL[308] WL[307] WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300]
+WL[299] WL[298] WL[297] WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] WL[290]
+WL[289] WL[288] WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] WL[281] WL[280]
+WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273] WL[272] WL[271] WL[270]
+WL[269] WL[268] WL[267] WL[266] WL[265] WL[264] WL[263] WL[262] WL[261] WL[260]
+WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_UP
XI14 UBL[3] UBL[2] UBLX[3] UBLX[2] RWLU[0] RWLU[1] VDD VSS WL[511] WL[510]
+WL[509] WL[508] WL[507] WL[506] WL[505] WL[504] WL[503] WL[502] WL[501] WL[500]
+WL[499] WL[498] WL[497] WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] WL[490]
+WL[489] WL[488] WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480]
+WL[479] WL[478] WL[477] WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] WL[470]
+WL[469] WL[468] WL[467] WL[466] WL[465] WL[464] WL[463] WL[462] WL[461] WL[460]
+WL[459] WL[458] WL[457] WL[456] WL[455] WL[454] WL[453] WL[452] WL[451] WL[450]
+WL[449] WL[448] WL[447] WL[446] WL[445] WL[444] WL[443] WL[442] WL[441] WL[440]
+WL[439] WL[438] WL[437] WL[436] WL[435] WL[434] WL[433] WL[432] WL[431] WL[430]
+WL[429] WL[428] WL[427] WL[426] WL[425] WL[424] WL[423] WL[422] WL[421] WL[420]
+WL[419] WL[418] WL[417] WL[416] WL[415] WL[414] WL[413] WL[412] WL[411] WL[410]
+WL[409] WL[408] WL[407] WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] WL[400]
+WL[399] WL[398] WL[397] WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390]
+WL[389] WL[388] WL[387] WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] WL[380]
+WL[379] WL[378] WL[377] WL[376] WL[375] WL[374] WL[373] WL[372] WL[371] WL[370]
+WL[369] WL[368] WL[367] WL[366] WL[365] WL[364] WL[363] WL[362] WL[361] WL[360]
+WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] WL[353] WL[352] WL[351] WL[350]
+WL[349] WL[348] WL[347] WL[346] WL[345] WL[344] WL[343] WL[342] WL[341] WL[340]
+WL[339] WL[338] WL[337] WL[336] WL[335] WL[334] WL[333] WL[332] WL[331] WL[330]
+WL[329] WL[328] WL[327] WL[326] WL[325] WL[324] WL[323] WL[322] WL[321] WL[320]
+WL[319] WL[318] WL[317] WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] WL[310]
+WL[309] WL[308] WL[307] WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300]
+WL[299] WL[298] WL[297] WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] WL[290]
+WL[289] WL[288] WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] WL[281] WL[280]
+WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273] WL[272] WL[271] WL[270]
+WL[269] WL[268] WL[267] WL[266] WL[265] WL[264] WL[263] WL[262] WL[261] WL[260]
+WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_UP
XI15 UBL[1] UBL[0] UBLX[1] UBLX[0] RWLU[0] RWLU[1] VDD VSS WL[511] WL[510]
+WL[509] WL[508] WL[507] WL[506] WL[505] WL[504] WL[503] WL[502] WL[501] WL[500]
+WL[499] WL[498] WL[497] WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] WL[490]
+WL[489] WL[488] WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480]
+WL[479] WL[478] WL[477] WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] WL[470]
+WL[469] WL[468] WL[467] WL[466] WL[465] WL[464] WL[463] WL[462] WL[461] WL[460]
+WL[459] WL[458] WL[457] WL[456] WL[455] WL[454] WL[453] WL[452] WL[451] WL[450]
+WL[449] WL[448] WL[447] WL[446] WL[445] WL[444] WL[443] WL[442] WL[441] WL[440]
+WL[439] WL[438] WL[437] WL[436] WL[435] WL[434] WL[433] WL[432] WL[431] WL[430]
+WL[429] WL[428] WL[427] WL[426] WL[425] WL[424] WL[423] WL[422] WL[421] WL[420]
+WL[419] WL[418] WL[417] WL[416] WL[415] WL[414] WL[413] WL[412] WL[411] WL[410]
+WL[409] WL[408] WL[407] WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] WL[400]
+WL[399] WL[398] WL[397] WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390]
+WL[389] WL[388] WL[387] WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] WL[380]
+WL[379] WL[378] WL[377] WL[376] WL[375] WL[374] WL[373] WL[372] WL[371] WL[370]
+WL[369] WL[368] WL[367] WL[366] WL[365] WL[364] WL[363] WL[362] WL[361] WL[360]
+WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] WL[353] WL[352] WL[351] WL[350]
+WL[349] WL[348] WL[347] WL[346] WL[345] WL[344] WL[343] WL[342] WL[341] WL[340]
+WL[339] WL[338] WL[337] WL[336] WL[335] WL[334] WL[333] WL[332] WL[331] WL[330]
+WL[329] WL[328] WL[327] WL[326] WL[325] WL[324] WL[323] WL[322] WL[321] WL[320]
+WL[319] WL[318] WL[317] WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] WL[310]
+WL[309] WL[308] WL[307] WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300]
+WL[299] WL[298] WL[297] WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] WL[290]
+WL[289] WL[288] WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] WL[281] WL[280]
+WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273] WL[272] WL[271] WL[270]
+WL[269] WL[268] WL[267] WL[266] WL[265] WL[264] WL[263] WL[262] WL[261] WL[260]
+WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_UP
XI16 DCTRCLK DCTRCLKX D[0] Q[0] LBL[15] LBL[14] LBL[13] LBL[12] LBL[11] LBL[10]
+LBL[9] LBL[8] LBL[7] LBL[6] LBL[5] LBL[4] LBL[3] LBL[2] LBL[1] LBL[0]
+LBLX[15] LBLX[14] LBLX[13] LBLX[12] LBLX[11] LBLX[10] LBLX[9] LBLX[8] LBLX[7] LBLX[6]
+LBLX[5] LBLX[4] LBLX[3] LBLX[2] LBLX[1] LBLX[0] SACK1 SACK4 UBL[15] UBL[14]
+UBL[13] UBL[12] UBL[11] UBL[10] UBL[9] UBL[8] UBL[7] UBL[6] UBL[5] UBL[4]
+UBL[3] UBL[2] UBL[1] UBL[0] UBLX[15] UBLX[14] UBLX[13] UBLX[12] UBLX[11] UBLX[10]
+UBLX[9] UBLX[8] UBLX[7] UBLX[6] UBLX[5] UBLX[4] UBLX[3] UBLX[2] UBLX[1] UBLX[0]
+VDD VSS WE YAX YX[7] YX[6] YX[5] YX[4] YX[3] YX[2]
+YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_YMX16SAWR
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP_EDGE256_UP
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP_EDGE256_UP RWL0 RWL1 VDD VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250]
+WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240]
+WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230]
+WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220]
+WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210]
+WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200]
+WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] WL[190]
+WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180]
+WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170]
+WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160]
+WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150]
+WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140]
+WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130]
+WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120]
+WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110]
+WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100]
+WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90]
+WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80]
+WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70]
+WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60]
+WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50]
+WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40]
+WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30]
+WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20]
+WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10]
+WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XI0 RWL0 RWL1 VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_PCAP_EDGE66B_RED
XI1 VDD VSS WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120]
+WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110]
+WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100]
+WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90]
+WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80]
+WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70]
+WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] S55NLLGSPH_X512Y16D32_PCAP_EDGE64A
XI2 VDD VSS WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184]
+WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174]
+WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164]
+WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154]
+WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144]
+WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134]
+WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] S55NLLGSPH_X512Y16D32_PCAP_EDGE64B
XI3 VDD VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248]
+WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238]
+WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228]
+WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218]
+WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208]
+WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198]
+WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] S55NLLGSPH_X512Y16D32_PCAP_EDGE64A
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_ARRAY_X512Y16D16_LEFT
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_ARRAY_X512Y16D16_LEFT D[15] D[14] D[13] D[12] D[11] D[10] D[9] D[8] D[7] D[6]
+D[5] D[4] D[3] D[2] D[1] D[0] DCTRCLK DCTRCLKX Q[15] Q[14]
+Q[13] Q[12] Q[11] Q[10] Q[9] Q[8] Q[7] Q[6] Q[5] Q[4]
+Q[3] Q[2] Q[1] Q[0] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX
XI0 RWLL[0] RWLL[1] STWL VDD VSS WL[255] WL[254] WL[253] WL[252] WL[251]
+WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241]
+WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231]
+WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221]
+WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211]
+WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201]
+WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191]
+WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181]
+WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171]
+WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161]
+WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151]
+WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141]
+WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131]
+WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121]
+WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111]
+WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101]
+WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91]
+WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81]
+WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71]
+WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61]
+WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51]
+WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41]
+WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31]
+WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21]
+WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11]
+WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1]
+WL[0] S55NLLGSPH_X512Y16D32_PCAP_EDGE256_DOWN
XI1 RWLL[0] RWLL[1] STWL VDD VSS WL[255] WL[254] WL[253] WL[252] WL[251]
+WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241]
+WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231]
+WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221]
+WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211]
+WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201]
+WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191]
+WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181]
+WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171]
+WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161]
+WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151]
+WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141]
+WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131]
+WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121]
+WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111]
+WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101]
+WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91]
+WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81]
+WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71]
+WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61]
+WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51]
+WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41]
+WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31]
+WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21]
+WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11]
+WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1]
+WL[0] S55NLLGSPH_X512Y16D32_PCAP_EDGE256_DOWN
XI2 D[0] DCTRCLK DCTRCLKX Q[0] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI3 D[1] DCTRCLK DCTRCLKX Q[1] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI4 D[2] DCTRCLK DCTRCLKX Q[2] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI5 D[3] DCTRCLK DCTRCLKX Q[3] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI6 D[4] DCTRCLK DCTRCLKX Q[4] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI7 D[5] DCTRCLK DCTRCLKX Q[5] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI8 D[6] DCTRCLK DCTRCLKX Q[6] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI9 D[7] DCTRCLK DCTRCLKX Q[7] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI10 D[8] DCTRCLK DCTRCLKX Q[8] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI11 D[9] DCTRCLK DCTRCLKX Q[9] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI12 D[10] DCTRCLK DCTRCLKX Q[10] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI13 D[11] DCTRCLK DCTRCLKX Q[11] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI14 D[12] DCTRCLK DCTRCLKX Q[12] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI15 D[13] DCTRCLK DCTRCLKX Q[13] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI16 D[14] DCTRCLK DCTRCLKX Q[14] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI17 D[15] DCTRCLK DCTRCLKX Q[15] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI18 RWLU[0] RWLU[1] VDD VSS WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_PCAP_EDGE256_UP
XI19 RWLU[0] RWLU[1] VDD VSS WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_PCAP_EDGE256_UP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP4A_ST
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP4A_ST BL VDD VSS WL[3] WL[2] WL[1] WL[0]
XI5 NET30 BL VDD VSS WL[3] S55NLLGSPH_X512Y16D32_PCAP
XI4 NET30 BL VDD VSS WL[2] S55NLLGSPH_X512Y16D32_PCAP
XI3 NET40 BL VDD VSS WL[1] S55NLLGSPH_X512Y16D32_PCAP
XI2 NET40 BL VDD VSS WL[0] S55NLLGSPH_X512Y16D32_PCAP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP64_ST
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP64_ST BL VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57]
+WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47]
+WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37]
+WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27]
+WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17]
+WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7]
+WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XI0 BL VDD VSS WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_PCAP4A_ST
XI1 BL VDD VSS WL[7] WL[6] WL[5] WL[4] S55NLLGSPH_X512Y16D32_PCAP4A_ST
XI2 BL VDD VSS WL[11] WL[10] WL[9] WL[8] S55NLLGSPH_X512Y16D32_PCAP4A_ST
XI3 BL VDD VSS WL[15] WL[14] WL[13] WL[12] S55NLLGSPH_X512Y16D32_PCAP4A_ST
XI4 BL VDD VSS WL[19] WL[18] WL[17] WL[16] S55NLLGSPH_X512Y16D32_PCAP4A_ST
XI5 BL VDD VSS WL[23] WL[22] WL[21] WL[20] S55NLLGSPH_X512Y16D32_PCAP4A_ST
XI6 BL VDD VSS WL[27] WL[26] WL[25] WL[24] S55NLLGSPH_X512Y16D32_PCAP4A_ST
XI7 BL VDD VSS WL[31] WL[30] WL[29] WL[28] S55NLLGSPH_X512Y16D32_PCAP4A_ST
XI8 BL VDD VSS WL[35] WL[34] WL[33] WL[32] S55NLLGSPH_X512Y16D32_PCAP4A_ST
XI9 BL VDD VSS WL[39] WL[38] WL[37] WL[36] S55NLLGSPH_X512Y16D32_PCAP4A_ST
XI10 BL VDD VSS WL[43] WL[42] WL[41] WL[40] S55NLLGSPH_X512Y16D32_PCAP4A_ST
XI11 BL VDD VSS WL[47] WL[46] WL[45] WL[44] S55NLLGSPH_X512Y16D32_PCAP4A_ST
XI12 BL VDD VSS WL[51] WL[50] WL[49] WL[48] S55NLLGSPH_X512Y16D32_PCAP4A_ST
XI13 BL VDD VSS WL[55] WL[54] WL[53] WL[52] S55NLLGSPH_X512Y16D32_PCAP4A_ST
XI14 BL VDD VSS WL[59] WL[58] WL[57] WL[56] S55NLLGSPH_X512Y16D32_PCAP4A_ST
XI15 BL VDD VSS WL[63] WL[62] WL[61] WL[60] S55NLLGSPH_X512Y16D32_PCAP4A_ST
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP_EDGE66A_ST_RED
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP_EDGE66A_ST_RED BL RWL0 RWL1 VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59]
+WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49]
+WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39]
+WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29]
+WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19]
+WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9]
+WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XI0 BL VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI1 BL VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57]
+WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47]
+WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37]
+WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27]
+WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17]
+WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7]
+WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_PCAP64_ST
XI2 NET43 BL VDD VSS RWL0 S55NLLGSPH_X512Y16D32_PCAP
XI3 NET43 BL VDD VSS RWL1 S55NLLGSPH_X512Y16D32_PCAP
XI4 BL VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP4B_ST
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP4B_ST BL BX0 BX1 VDD VSS WL[3] WL[2] WL[1] WL[0]
XI5 BX1 BL VDD VSS WL[3] S55NLLGSPH_X512Y16D32_PCAP
XI4 NET37 BL VDD VSS WL[2] S55NLLGSPH_X512Y16D32_PCAP
XI3 NET37 BL VDD VSS WL[1] S55NLLGSPH_X512Y16D32_PCAP
XI2 BX0 BL VDD VSS WL[0] S55NLLGSPH_X512Y16D32_PCAP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP64B_ST
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP64B_ST BL BX0 BX1 VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59]
+WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49]
+WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39]
+WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29]
+WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19]
+WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9]
+WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XI0 BL NET31 NET61 VDD VSS WL[7] WL[6] WL[5] WL[4] S55NLLGSPH_X512Y16D32_PCAP4B_ST
XI1 BL BX0 NET31 VDD VSS WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_PCAP4B_ST
XI2 BL NET01 NET32 VDD VSS WL[11] WL[10] WL[9] WL[8] S55NLLGSPH_X512Y16D32_PCAP4B_ST
XI3 BL NET32 NET61 VDD VSS WL[15] WL[14] WL[13] WL[12] S55NLLGSPH_X512Y16D32_PCAP4B_ST
XI4 BL NET33 NET62 VDD VSS WL[23] WL[22] WL[21] WL[20] S55NLLGSPH_X512Y16D32_PCAP4B_ST
XI5 BL NET01 NET33 VDD VSS WL[19] WL[18] WL[17] WL[16] S55NLLGSPH_X512Y16D32_PCAP4B_ST
XI6 BL NET02 NET34 VDD VSS WL[27] WL[26] WL[25] WL[24] S55NLLGSPH_X512Y16D32_PCAP4B_ST
XI7 BL NET34 NET62 VDD VSS WL[31] WL[30] WL[29] WL[28] S55NLLGSPH_X512Y16D32_PCAP4B_ST
XI8 BL NET35 NET63 VDD VSS WL[39] WL[38] WL[37] WL[36] S55NLLGSPH_X512Y16D32_PCAP4B_ST
XI9 BL NET02 NET35 VDD VSS WL[35] WL[34] WL[33] WL[32] S55NLLGSPH_X512Y16D32_PCAP4B_ST
XI10 BL NET03 NET36 VDD VSS WL[43] WL[42] WL[41] WL[40] S55NLLGSPH_X512Y16D32_PCAP4B_ST
XI11 BL NET36 NET63 VDD VSS WL[47] WL[46] WL[45] WL[44] S55NLLGSPH_X512Y16D32_PCAP4B_ST
XI12 BL NET37 NET64 VDD VSS WL[55] WL[54] WL[53] WL[52] S55NLLGSPH_X512Y16D32_PCAP4B_ST
XI13 BL NET03 NET37 VDD VSS WL[51] WL[50] WL[49] WL[48] S55NLLGSPH_X512Y16D32_PCAP4B_ST
XI14 BL BX1 NET38 VDD VSS WL[59] WL[58] WL[57] WL[56] S55NLLGSPH_X512Y16D32_PCAP4B_ST
XI15 BL NET38 NET64 VDD VSS WL[63] WL[62] WL[61] WL[60] S55NLLGSPH_X512Y16D32_PCAP4B_ST
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP_EDGE64B_ST
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP_EDGE64B_ST BL VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57]
+WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47]
+WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37]
+WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27]
+WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17]
+WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7]
+WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XI0 NET28 VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI1 BL NET28 NET024 VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59]
+WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49]
+WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39]
+WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29]
+WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19]
+WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9]
+WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_PCAP64B_ST
XI2 NET024 VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP_EDGE64A_ST
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP_EDGE64A_ST BL VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57]
+WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47]
+WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37]
+WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27]
+WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17]
+WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7]
+WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XI0 BL VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI1 BL VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57]
+WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47]
+WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37]
+WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27]
+WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17]
+WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7]
+WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_PCAP64_ST
XI2 BL VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP4B_ST_RDWL
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP4B_ST_RDWL BX0 BX1 VDD VSS WL[0] WL[1] WL[2] WL[3]
XI5 BX1 NET031 VDD VSS WL[3] S55NLLGSPH_X512Y16D32_PCAP
XI4 NET37 NET031 VDD VSS WL[2] S55NLLGSPH_X512Y16D32_PCAP
XI3 NET37 NET041 VDD VSS WL[1] S55NLLGSPH_X512Y16D32_PCAP
XI2 BX0 NET041 VDD VSS WL[0] S55NLLGSPH_X512Y16D32_PCAP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP_EDGE68B_ST_TOP
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP_EDGE68B_ST_TOP BL RDWL VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XI0 NET28 VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI1 BL NET28 NET024 VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59]
+WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49]
+WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39]
+WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29]
+WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19]
+WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9]
+WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_PCAP64B_ST
XI2 NET024 NET39 VDD VSS VSS RDWL RDWL VSS S55NLLGSPH_X512Y16D32_PCAP4B_ST_RDWL
XI3 NET39 VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PCAP_EDGE256_ST
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PCAP_EDGE256_ST BL RWL0 RWL1 STWL VDD VSS WL[255] WL[254] WL[253] WL[252]
+WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243] WL[242]
+WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233] WL[232]
+WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223] WL[222]
+WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213] WL[212]
+WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] WL[202]
+WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192]
+WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183] WL[182]
+WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173] WL[172]
+WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163] WL[162]
+WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153] WL[152]
+WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143] WL[142]
+WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133] WL[132]
+WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123] WL[122]
+WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] WL[112]
+WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102]
+WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92]
+WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82]
+WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72]
+WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63] WL[62]
+WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52]
+WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42]
+WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32]
+WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22]
+WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12]
+WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2]
+WL[1] WL[0]
XI0 BL RWL0 RWL1 VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59]
+WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49]
+WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39]
+WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29]
+WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19]
+WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9]
+WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_PCAP_EDGE66A_ST_RED
XI1 BL VDD VSS WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121]
+WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111]
+WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101]
+WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91]
+WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81]
+WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71]
+WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] S55NLLGSPH_X512Y16D32_PCAP_EDGE64B_ST
XI2 BL VDD VSS WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] S55NLLGSPH_X512Y16D32_PCAP_EDGE64A_ST
XI3 BL STWL VDD VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250]
+WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240]
+WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230]
+WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220]
+WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210]
+WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200]
+WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] S55NLLGSPH_X512Y16D32_PCAP_EDGE68B_ST_TOP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525_MD
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525_MD B BX VDD VSS WL0 WL1
MM2 BX WL0 BCN VSS STNPGHVT W=85.000N L=75.00N M=1
MM3 B WL1 BC VSS STNPGHVT W=85.000N L=75.00N M=1
MM0 BCN BC VSS VSS STNPDHVT W=135.00N L=65.00N M=1
MM1 BC BCN VSS VSS STNPDHVT W=135.00N L=65.00N M=1
MM5 BCN BC VDD VDD STPLHVT W=85.000N L=65.00N M=1
MM6 BC BCN VDD VDD STPLHVT W=85.000N L=65.00N M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_BITCELL_RDWL2B_MD
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_BITCELL_RDWL2B_MD BLL[1] BLL[0] BLU[1] BLU[0] VDD VSS WL0 WL1 WL2 WL3
XI2 NET034 NET028 VDD VSS WL2 VSS S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525_MD
XI1 NET034 NET043 VDD VSS WL1 VSS S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525_MD
XI7 BLL[1] NET018 VDD VSS WL3 S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525
XI4 NET024 NET018 VDD VSS WL2 S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525
XI9 BLL[0] NET028 VDD VSS VSS S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525
XI8 BLU[0] NET043 VDD VSS VSS S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525
XI5 BLU[1] NET11 VDD VSS WL0 S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525
XI6 NET024 NET11 VDD VSS WL1 S55NLLGSPH_X512Y16D32_BITCELL_HSSPH_HVT525
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_BITCELL68X2B_TOP_MD
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_BITCELL68X2B_TOP_MD BL[1] BL[0] BLX[1] BLX[0] RDWL VDD VSS WL[63] WL[62] WL[61]
+WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51]
+WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41]
+WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31]
+WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21]
+WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11]
+WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1]
+WL[0]
XI0 NET47[0] NET47[1] BL[1] BL[0] VDD VSS VSS RDWL RDWL VSS S55NLLGSPH_X512Y16D32_BITCELL_RDWL2B_MD
XI1 NET47[0] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI2 NET47[1] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI3 BL[1] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI4 BL[0] VDD VSS S55NLLGSPH_X512Y16D32_BLSTRAP1
XI5 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI6 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[3] WL[2] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI7 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[5] WL[4] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI8 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[7] WL[6] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI9 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[9] WL[8] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI10 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[11] WL[10] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI11 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[13] WL[12] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI12 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[15] WL[14] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI13 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[17] WL[16] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI14 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[19] WL[18] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI15 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[21] WL[20] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI16 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[23] WL[22] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI17 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[25] WL[24] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI18 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[27] WL[26] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI19 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[29] WL[28] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI20 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[31] WL[30] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI21 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[33] WL[32] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI22 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[35] WL[34] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI23 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[37] WL[36] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI24 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[39] WL[38] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI25 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[41] WL[40] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI26 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[43] WL[42] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI27 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[45] WL[44] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI28 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[47] WL[46] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI29 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[49] WL[48] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI30 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[51] WL[50] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI31 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[53] WL[52] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI32 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[55] WL[54] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI33 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[57] WL[56] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI34 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[59] WL[58] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI35 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[61] WL[60] S55NLLGSPH_X512Y16D32_BITCELL2X2
XI36 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[63] WL[62] S55NLLGSPH_X512Y16D32_BITCELL2X2
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN_MD
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN_MD BL[1] BL[0] BLX[1] BLX[0] RDWL RWL[0] RWL[1] VDD VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0]
XI0 BL[1] BL[0] BLX[1] BLX[0] RWL[0] RWL[1] VDD VSS WL[63] WL[62]
+WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52]
+WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42]
+WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32]
+WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22]
+WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12]
+WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2]
+WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL66X2A_RED
XI1 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[127] WL[126] WL[125] WL[124]
+WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114]
+WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104]
+WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94]
+WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84]
+WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74]
+WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] S55NLLGSPH_X512Y16D32_BITCELL64X2B
XI2 BL[1] BL[0] BLX[1] BLX[0] VDD VSS WL[191] WL[190] WL[189] WL[188]
+WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178]
+WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168]
+WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158]
+WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148]
+WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138]
+WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] S55NLLGSPH_X512Y16D32_BITCELL64X2A
XI3 BL[1] BL[0] BLX[1] BLX[0] RDWL VDD VSS WL[255] WL[254] WL[253]
+WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243]
+WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223]
+WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213]
+WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203]
+WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] S55NLLGSPH_X512Y16D32_BITCELL68X2B_TOP_MD
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_Y16_X512_D1_MD
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_Y16_X512_D1_MD D[0] DCTRCLK DCTRCLKX Q[0] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX
XI0 LBL[15] LBL[14] LBLX[15] LBLX[14] STWL RWLL[0] RWLL[1] VDD VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN
XI1 LBL[13] LBL[12] LBLX[13] LBLX[12] STWL RWLL[0] RWLL[1] VDD VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN
XI2 LBL[11] LBL[10] LBLX[11] LBLX[10] STWL RWLL[0] RWLL[1] VDD VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN
XI3 LBL[9] LBL[8] LBLX[9] LBLX[8] STWL RWLL[0] RWLL[1] VDD VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN
XI4 LBL[7] LBL[6] LBLX[7] LBLX[6] STWL RWLL[0] RWLL[1] VDD VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN
XI5 LBL[5] LBL[4] LBLX[5] LBLX[4] STWL RWLL[0] RWLL[1] VDD VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN
XI6 LBL[3] LBL[2] LBLX[3] LBLX[2] STWL RWLL[0] RWLL[1] VDD VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN
XI7 LBL[1] LBL[0] LBLX[1] LBLX[0] STWL RWLL[0] RWLL[1] VDD VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_DOWN_MD
XI8 UBL[15] UBL[14] UBLX[15] UBLX[14] RWLU[0] RWLU[1] VDD VSS WL[511] WL[510]
+WL[509] WL[508] WL[507] WL[506] WL[505] WL[504] WL[503] WL[502] WL[501] WL[500]
+WL[499] WL[498] WL[497] WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] WL[490]
+WL[489] WL[488] WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480]
+WL[479] WL[478] WL[477] WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] WL[470]
+WL[469] WL[468] WL[467] WL[466] WL[465] WL[464] WL[463] WL[462] WL[461] WL[460]
+WL[459] WL[458] WL[457] WL[456] WL[455] WL[454] WL[453] WL[452] WL[451] WL[450]
+WL[449] WL[448] WL[447] WL[446] WL[445] WL[444] WL[443] WL[442] WL[441] WL[440]
+WL[439] WL[438] WL[437] WL[436] WL[435] WL[434] WL[433] WL[432] WL[431] WL[430]
+WL[429] WL[428] WL[427] WL[426] WL[425] WL[424] WL[423] WL[422] WL[421] WL[420]
+WL[419] WL[418] WL[417] WL[416] WL[415] WL[414] WL[413] WL[412] WL[411] WL[410]
+WL[409] WL[408] WL[407] WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] WL[400]
+WL[399] WL[398] WL[397] WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390]
+WL[389] WL[388] WL[387] WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] WL[380]
+WL[379] WL[378] WL[377] WL[376] WL[375] WL[374] WL[373] WL[372] WL[371] WL[370]
+WL[369] WL[368] WL[367] WL[366] WL[365] WL[364] WL[363] WL[362] WL[361] WL[360]
+WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] WL[353] WL[352] WL[351] WL[350]
+WL[349] WL[348] WL[347] WL[346] WL[345] WL[344] WL[343] WL[342] WL[341] WL[340]
+WL[339] WL[338] WL[337] WL[336] WL[335] WL[334] WL[333] WL[332] WL[331] WL[330]
+WL[329] WL[328] WL[327] WL[326] WL[325] WL[324] WL[323] WL[322] WL[321] WL[320]
+WL[319] WL[318] WL[317] WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] WL[310]
+WL[309] WL[308] WL[307] WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300]
+WL[299] WL[298] WL[297] WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] WL[290]
+WL[289] WL[288] WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] WL[281] WL[280]
+WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273] WL[272] WL[271] WL[270]
+WL[269] WL[268] WL[267] WL[266] WL[265] WL[264] WL[263] WL[262] WL[261] WL[260]
+WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_UP
XI9 UBL[13] UBL[12] UBLX[13] UBLX[12] RWLU[0] RWLU[1] VDD VSS WL[511] WL[510]
+WL[509] WL[508] WL[507] WL[506] WL[505] WL[504] WL[503] WL[502] WL[501] WL[500]
+WL[499] WL[498] WL[497] WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] WL[490]
+WL[489] WL[488] WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480]
+WL[479] WL[478] WL[477] WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] WL[470]
+WL[469] WL[468] WL[467] WL[466] WL[465] WL[464] WL[463] WL[462] WL[461] WL[460]
+WL[459] WL[458] WL[457] WL[456] WL[455] WL[454] WL[453] WL[452] WL[451] WL[450]
+WL[449] WL[448] WL[447] WL[446] WL[445] WL[444] WL[443] WL[442] WL[441] WL[440]
+WL[439] WL[438] WL[437] WL[436] WL[435] WL[434] WL[433] WL[432] WL[431] WL[430]
+WL[429] WL[428] WL[427] WL[426] WL[425] WL[424] WL[423] WL[422] WL[421] WL[420]
+WL[419] WL[418] WL[417] WL[416] WL[415] WL[414] WL[413] WL[412] WL[411] WL[410]
+WL[409] WL[408] WL[407] WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] WL[400]
+WL[399] WL[398] WL[397] WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390]
+WL[389] WL[388] WL[387] WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] WL[380]
+WL[379] WL[378] WL[377] WL[376] WL[375] WL[374] WL[373] WL[372] WL[371] WL[370]
+WL[369] WL[368] WL[367] WL[366] WL[365] WL[364] WL[363] WL[362] WL[361] WL[360]
+WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] WL[353] WL[352] WL[351] WL[350]
+WL[349] WL[348] WL[347] WL[346] WL[345] WL[344] WL[343] WL[342] WL[341] WL[340]
+WL[339] WL[338] WL[337] WL[336] WL[335] WL[334] WL[333] WL[332] WL[331] WL[330]
+WL[329] WL[328] WL[327] WL[326] WL[325] WL[324] WL[323] WL[322] WL[321] WL[320]
+WL[319] WL[318] WL[317] WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] WL[310]
+WL[309] WL[308] WL[307] WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300]
+WL[299] WL[298] WL[297] WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] WL[290]
+WL[289] WL[288] WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] WL[281] WL[280]
+WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273] WL[272] WL[271] WL[270]
+WL[269] WL[268] WL[267] WL[266] WL[265] WL[264] WL[263] WL[262] WL[261] WL[260]
+WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_UP
XI10 UBL[11] UBL[10] UBLX[11] UBLX[10] RWLU[0] RWLU[1] VDD VSS WL[511] WL[510]
+WL[509] WL[508] WL[507] WL[506] WL[505] WL[504] WL[503] WL[502] WL[501] WL[500]
+WL[499] WL[498] WL[497] WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] WL[490]
+WL[489] WL[488] WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480]
+WL[479] WL[478] WL[477] WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] WL[470]
+WL[469] WL[468] WL[467] WL[466] WL[465] WL[464] WL[463] WL[462] WL[461] WL[460]
+WL[459] WL[458] WL[457] WL[456] WL[455] WL[454] WL[453] WL[452] WL[451] WL[450]
+WL[449] WL[448] WL[447] WL[446] WL[445] WL[444] WL[443] WL[442] WL[441] WL[440]
+WL[439] WL[438] WL[437] WL[436] WL[435] WL[434] WL[433] WL[432] WL[431] WL[430]
+WL[429] WL[428] WL[427] WL[426] WL[425] WL[424] WL[423] WL[422] WL[421] WL[420]
+WL[419] WL[418] WL[417] WL[416] WL[415] WL[414] WL[413] WL[412] WL[411] WL[410]
+WL[409] WL[408] WL[407] WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] WL[400]
+WL[399] WL[398] WL[397] WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390]
+WL[389] WL[388] WL[387] WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] WL[380]
+WL[379] WL[378] WL[377] WL[376] WL[375] WL[374] WL[373] WL[372] WL[371] WL[370]
+WL[369] WL[368] WL[367] WL[366] WL[365] WL[364] WL[363] WL[362] WL[361] WL[360]
+WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] WL[353] WL[352] WL[351] WL[350]
+WL[349] WL[348] WL[347] WL[346] WL[345] WL[344] WL[343] WL[342] WL[341] WL[340]
+WL[339] WL[338] WL[337] WL[336] WL[335] WL[334] WL[333] WL[332] WL[331] WL[330]
+WL[329] WL[328] WL[327] WL[326] WL[325] WL[324] WL[323] WL[322] WL[321] WL[320]
+WL[319] WL[318] WL[317] WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] WL[310]
+WL[309] WL[308] WL[307] WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300]
+WL[299] WL[298] WL[297] WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] WL[290]
+WL[289] WL[288] WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] WL[281] WL[280]
+WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273] WL[272] WL[271] WL[270]
+WL[269] WL[268] WL[267] WL[266] WL[265] WL[264] WL[263] WL[262] WL[261] WL[260]
+WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_UP
XI11 UBL[9] UBL[8] UBLX[9] UBLX[8] RWLU[0] RWLU[1] VDD VSS WL[511] WL[510]
+WL[509] WL[508] WL[507] WL[506] WL[505] WL[504] WL[503] WL[502] WL[501] WL[500]
+WL[499] WL[498] WL[497] WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] WL[490]
+WL[489] WL[488] WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480]
+WL[479] WL[478] WL[477] WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] WL[470]
+WL[469] WL[468] WL[467] WL[466] WL[465] WL[464] WL[463] WL[462] WL[461] WL[460]
+WL[459] WL[458] WL[457] WL[456] WL[455] WL[454] WL[453] WL[452] WL[451] WL[450]
+WL[449] WL[448] WL[447] WL[446] WL[445] WL[444] WL[443] WL[442] WL[441] WL[440]
+WL[439] WL[438] WL[437] WL[436] WL[435] WL[434] WL[433] WL[432] WL[431] WL[430]
+WL[429] WL[428] WL[427] WL[426] WL[425] WL[424] WL[423] WL[422] WL[421] WL[420]
+WL[419] WL[418] WL[417] WL[416] WL[415] WL[414] WL[413] WL[412] WL[411] WL[410]
+WL[409] WL[408] WL[407] WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] WL[400]
+WL[399] WL[398] WL[397] WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390]
+WL[389] WL[388] WL[387] WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] WL[380]
+WL[379] WL[378] WL[377] WL[376] WL[375] WL[374] WL[373] WL[372] WL[371] WL[370]
+WL[369] WL[368] WL[367] WL[366] WL[365] WL[364] WL[363] WL[362] WL[361] WL[360]
+WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] WL[353] WL[352] WL[351] WL[350]
+WL[349] WL[348] WL[347] WL[346] WL[345] WL[344] WL[343] WL[342] WL[341] WL[340]
+WL[339] WL[338] WL[337] WL[336] WL[335] WL[334] WL[333] WL[332] WL[331] WL[330]
+WL[329] WL[328] WL[327] WL[326] WL[325] WL[324] WL[323] WL[322] WL[321] WL[320]
+WL[319] WL[318] WL[317] WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] WL[310]
+WL[309] WL[308] WL[307] WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300]
+WL[299] WL[298] WL[297] WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] WL[290]
+WL[289] WL[288] WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] WL[281] WL[280]
+WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273] WL[272] WL[271] WL[270]
+WL[269] WL[268] WL[267] WL[266] WL[265] WL[264] WL[263] WL[262] WL[261] WL[260]
+WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_UP
XI12 UBL[7] UBL[6] UBLX[7] UBLX[6] RWLU[0] RWLU[1] VDD VSS WL[511] WL[510]
+WL[509] WL[508] WL[507] WL[506] WL[505] WL[504] WL[503] WL[502] WL[501] WL[500]
+WL[499] WL[498] WL[497] WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] WL[490]
+WL[489] WL[488] WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480]
+WL[479] WL[478] WL[477] WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] WL[470]
+WL[469] WL[468] WL[467] WL[466] WL[465] WL[464] WL[463] WL[462] WL[461] WL[460]
+WL[459] WL[458] WL[457] WL[456] WL[455] WL[454] WL[453] WL[452] WL[451] WL[450]
+WL[449] WL[448] WL[447] WL[446] WL[445] WL[444] WL[443] WL[442] WL[441] WL[440]
+WL[439] WL[438] WL[437] WL[436] WL[435] WL[434] WL[433] WL[432] WL[431] WL[430]
+WL[429] WL[428] WL[427] WL[426] WL[425] WL[424] WL[423] WL[422] WL[421] WL[420]
+WL[419] WL[418] WL[417] WL[416] WL[415] WL[414] WL[413] WL[412] WL[411] WL[410]
+WL[409] WL[408] WL[407] WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] WL[400]
+WL[399] WL[398] WL[397] WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390]
+WL[389] WL[388] WL[387] WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] WL[380]
+WL[379] WL[378] WL[377] WL[376] WL[375] WL[374] WL[373] WL[372] WL[371] WL[370]
+WL[369] WL[368] WL[367] WL[366] WL[365] WL[364] WL[363] WL[362] WL[361] WL[360]
+WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] WL[353] WL[352] WL[351] WL[350]
+WL[349] WL[348] WL[347] WL[346] WL[345] WL[344] WL[343] WL[342] WL[341] WL[340]
+WL[339] WL[338] WL[337] WL[336] WL[335] WL[334] WL[333] WL[332] WL[331] WL[330]
+WL[329] WL[328] WL[327] WL[326] WL[325] WL[324] WL[323] WL[322] WL[321] WL[320]
+WL[319] WL[318] WL[317] WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] WL[310]
+WL[309] WL[308] WL[307] WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300]
+WL[299] WL[298] WL[297] WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] WL[290]
+WL[289] WL[288] WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] WL[281] WL[280]
+WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273] WL[272] WL[271] WL[270]
+WL[269] WL[268] WL[267] WL[266] WL[265] WL[264] WL[263] WL[262] WL[261] WL[260]
+WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_UP
XI13 UBL[5] UBL[4] UBLX[5] UBLX[4] RWLU[0] RWLU[1] VDD VSS WL[511] WL[510]
+WL[509] WL[508] WL[507] WL[506] WL[505] WL[504] WL[503] WL[502] WL[501] WL[500]
+WL[499] WL[498] WL[497] WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] WL[490]
+WL[489] WL[488] WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480]
+WL[479] WL[478] WL[477] WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] WL[470]
+WL[469] WL[468] WL[467] WL[466] WL[465] WL[464] WL[463] WL[462] WL[461] WL[460]
+WL[459] WL[458] WL[457] WL[456] WL[455] WL[454] WL[453] WL[452] WL[451] WL[450]
+WL[449] WL[448] WL[447] WL[446] WL[445] WL[444] WL[443] WL[442] WL[441] WL[440]
+WL[439] WL[438] WL[437] WL[436] WL[435] WL[434] WL[433] WL[432] WL[431] WL[430]
+WL[429] WL[428] WL[427] WL[426] WL[425] WL[424] WL[423] WL[422] WL[421] WL[420]
+WL[419] WL[418] WL[417] WL[416] WL[415] WL[414] WL[413] WL[412] WL[411] WL[410]
+WL[409] WL[408] WL[407] WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] WL[400]
+WL[399] WL[398] WL[397] WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390]
+WL[389] WL[388] WL[387] WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] WL[380]
+WL[379] WL[378] WL[377] WL[376] WL[375] WL[374] WL[373] WL[372] WL[371] WL[370]
+WL[369] WL[368] WL[367] WL[366] WL[365] WL[364] WL[363] WL[362] WL[361] WL[360]
+WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] WL[353] WL[352] WL[351] WL[350]
+WL[349] WL[348] WL[347] WL[346] WL[345] WL[344] WL[343] WL[342] WL[341] WL[340]
+WL[339] WL[338] WL[337] WL[336] WL[335] WL[334] WL[333] WL[332] WL[331] WL[330]
+WL[329] WL[328] WL[327] WL[326] WL[325] WL[324] WL[323] WL[322] WL[321] WL[320]
+WL[319] WL[318] WL[317] WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] WL[310]
+WL[309] WL[308] WL[307] WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300]
+WL[299] WL[298] WL[297] WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] WL[290]
+WL[289] WL[288] WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] WL[281] WL[280]
+WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273] WL[272] WL[271] WL[270]
+WL[269] WL[268] WL[267] WL[266] WL[265] WL[264] WL[263] WL[262] WL[261] WL[260]
+WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_UP
XI14 UBL[3] UBL[2] UBLX[3] UBLX[2] RWLU[0] RWLU[1] VDD VSS WL[511] WL[510]
+WL[509] WL[508] WL[507] WL[506] WL[505] WL[504] WL[503] WL[502] WL[501] WL[500]
+WL[499] WL[498] WL[497] WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] WL[490]
+WL[489] WL[488] WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480]
+WL[479] WL[478] WL[477] WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] WL[470]
+WL[469] WL[468] WL[467] WL[466] WL[465] WL[464] WL[463] WL[462] WL[461] WL[460]
+WL[459] WL[458] WL[457] WL[456] WL[455] WL[454] WL[453] WL[452] WL[451] WL[450]
+WL[449] WL[448] WL[447] WL[446] WL[445] WL[444] WL[443] WL[442] WL[441] WL[440]
+WL[439] WL[438] WL[437] WL[436] WL[435] WL[434] WL[433] WL[432] WL[431] WL[430]
+WL[429] WL[428] WL[427] WL[426] WL[425] WL[424] WL[423] WL[422] WL[421] WL[420]
+WL[419] WL[418] WL[417] WL[416] WL[415] WL[414] WL[413] WL[412] WL[411] WL[410]
+WL[409] WL[408] WL[407] WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] WL[400]
+WL[399] WL[398] WL[397] WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390]
+WL[389] WL[388] WL[387] WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] WL[380]
+WL[379] WL[378] WL[377] WL[376] WL[375] WL[374] WL[373] WL[372] WL[371] WL[370]
+WL[369] WL[368] WL[367] WL[366] WL[365] WL[364] WL[363] WL[362] WL[361] WL[360]
+WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] WL[353] WL[352] WL[351] WL[350]
+WL[349] WL[348] WL[347] WL[346] WL[345] WL[344] WL[343] WL[342] WL[341] WL[340]
+WL[339] WL[338] WL[337] WL[336] WL[335] WL[334] WL[333] WL[332] WL[331] WL[330]
+WL[329] WL[328] WL[327] WL[326] WL[325] WL[324] WL[323] WL[322] WL[321] WL[320]
+WL[319] WL[318] WL[317] WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] WL[310]
+WL[309] WL[308] WL[307] WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300]
+WL[299] WL[298] WL[297] WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] WL[290]
+WL[289] WL[288] WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] WL[281] WL[280]
+WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273] WL[272] WL[271] WL[270]
+WL[269] WL[268] WL[267] WL[266] WL[265] WL[264] WL[263] WL[262] WL[261] WL[260]
+WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_UP
XI15 UBL[1] UBL[0] UBLX[1] UBLX[0] RWLU[0] RWLU[1] VDD VSS WL[511] WL[510]
+WL[509] WL[508] WL[507] WL[506] WL[505] WL[504] WL[503] WL[502] WL[501] WL[500]
+WL[499] WL[498] WL[497] WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] WL[490]
+WL[489] WL[488] WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480]
+WL[479] WL[478] WL[477] WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] WL[470]
+WL[469] WL[468] WL[467] WL[466] WL[465] WL[464] WL[463] WL[462] WL[461] WL[460]
+WL[459] WL[458] WL[457] WL[456] WL[455] WL[454] WL[453] WL[452] WL[451] WL[450]
+WL[449] WL[448] WL[447] WL[446] WL[445] WL[444] WL[443] WL[442] WL[441] WL[440]
+WL[439] WL[438] WL[437] WL[436] WL[435] WL[434] WL[433] WL[432] WL[431] WL[430]
+WL[429] WL[428] WL[427] WL[426] WL[425] WL[424] WL[423] WL[422] WL[421] WL[420]
+WL[419] WL[418] WL[417] WL[416] WL[415] WL[414] WL[413] WL[412] WL[411] WL[410]
+WL[409] WL[408] WL[407] WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] WL[400]
+WL[399] WL[398] WL[397] WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390]
+WL[389] WL[388] WL[387] WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] WL[380]
+WL[379] WL[378] WL[377] WL[376] WL[375] WL[374] WL[373] WL[372] WL[371] WL[370]
+WL[369] WL[368] WL[367] WL[366] WL[365] WL[364] WL[363] WL[362] WL[361] WL[360]
+WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] WL[353] WL[352] WL[351] WL[350]
+WL[349] WL[348] WL[347] WL[346] WL[345] WL[344] WL[343] WL[342] WL[341] WL[340]
+WL[339] WL[338] WL[337] WL[336] WL[335] WL[334] WL[333] WL[332] WL[331] WL[330]
+WL[329] WL[328] WL[327] WL[326] WL[325] WL[324] WL[323] WL[322] WL[321] WL[320]
+WL[319] WL[318] WL[317] WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] WL[310]
+WL[309] WL[308] WL[307] WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300]
+WL[299] WL[298] WL[297] WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] WL[290]
+WL[289] WL[288] WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] WL[281] WL[280]
+WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273] WL[272] WL[271] WL[270]
+WL[269] WL[268] WL[267] WL[266] WL[265] WL[264] WL[263] WL[262] WL[261] WL[260]
+WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_BITCELL256X2ABR_UP
XI16 DCTRCLK DCTRCLKX D[0] Q[0] LBL[15] LBL[14] LBL[13] LBL[12] LBL[11] LBL[10]
+LBL[9] LBL[8] LBL[7] LBL[6] LBL[5] LBL[4] LBL[3] LBL[2] LBL[1] LBL[0]
+LBLX[15] LBLX[14] LBLX[13] LBLX[12] LBLX[11] LBLX[10] LBLX[9] LBLX[8] LBLX[7] LBLX[6]
+LBLX[5] LBLX[4] LBLX[3] LBLX[2] LBLX[1] LBLX[0] SACK1 SACK4 UBL[15] UBL[14]
+UBL[13] UBL[12] UBL[11] UBL[10] UBL[9] UBL[8] UBL[7] UBL[6] UBL[5] UBL[4]
+UBL[3] UBL[2] UBL[1] UBL[0] UBLX[15] UBLX[14] UBLX[13] UBLX[12] UBLX[11] UBLX[10]
+UBLX[9] UBLX[8] UBLX[7] UBLX[6] UBLX[5] UBLX[4] UBLX[3] UBLX[2] UBLX[1] UBLX[0]
+VDD VSS WE YAX YX[7] YX[6] YX[5] YX[4] YX[3] YX[2]
+YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_YMX16SAWR
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_ARRAY_X512Y16D16_RIGHT
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_ARRAY_X512Y16D16_RIGHT D[15] D[14] D[13] D[12] D[11] D[10] D[9] D[8] D[7] D[6]
+D[5] D[4] D[3] D[2] D[1] D[0] DBL DCTRCLK DCTRCLKX Q[15]
+Q[14] Q[13] Q[12] Q[11] Q[10] Q[9] Q[8] Q[7] Q[6] Q[5]
+Q[4] Q[3] Q[2] Q[1] Q[0] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1
+SACK4 STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507]
+WL[506] WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497]
+WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487]
+WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477]
+WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467]
+WL[466] WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457]
+WL[456] WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447]
+WL[446] WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437]
+WL[436] WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427]
+WL[426] WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417]
+WL[416] WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407]
+WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397]
+WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387]
+WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377]
+WL[376] WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367]
+WL[366] WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357]
+WL[356] WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347]
+WL[346] WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337]
+WL[336] WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327]
+WL[326] WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317]
+WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307]
+WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297]
+WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287]
+WL[286] WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277]
+WL[276] WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267]
+WL[266] WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257]
+WL[256] WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247]
+WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237]
+WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227]
+WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217]
+WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207]
+WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197]
+WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187]
+WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177]
+WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167]
+WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157]
+WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147]
+WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137]
+WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127]
+WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117]
+WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107]
+WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97]
+WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87]
+WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77]
+WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67]
+WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57]
+WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47]
+WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37]
+WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27]
+WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17]
+WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7]
+WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6]
+YX[5] YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX
XI0 DBL RWLL[0] RWLL[1] STWL VDD VSS WL[255] WL[254] WL[253] WL[252]
+WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243] WL[242]
+WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233] WL[232]
+WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223] WL[222]
+WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213] WL[212]
+WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] WL[202]
+WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192]
+WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183] WL[182]
+WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173] WL[172]
+WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163] WL[162]
+WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153] WL[152]
+WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143] WL[142]
+WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133] WL[132]
+WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123] WL[122]
+WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] WL[112]
+WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102]
+WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92]
+WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82]
+WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72]
+WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63] WL[62]
+WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52]
+WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42]
+WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32]
+WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22]
+WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12]
+WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2]
+WL[1] WL[0] S55NLLGSPH_X512Y16D32_PCAP_EDGE256_ST
XI1 RWLL[0] RWLL[1] VSS VDD VSS WL[255] WL[254] WL[253] WL[252] WL[251]
+WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241]
+WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231]
+WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221]
+WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211]
+WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201]
+WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191]
+WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181]
+WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171]
+WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161]
+WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151]
+WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141]
+WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131]
+WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121]
+WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111]
+WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101]
+WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91]
+WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81]
+WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71]
+WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61]
+WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51]
+WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41]
+WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31]
+WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21]
+WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11]
+WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1]
+WL[0] S55NLLGSPH_X512Y16D32_PCAP_EDGE256_DOWN
XI2 D[0] DCTRCLK DCTRCLKX Q[0] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI3 D[1] DCTRCLK DCTRCLKX Q[1] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI4 D[2] DCTRCLK DCTRCLKX Q[2] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI5 D[3] DCTRCLK DCTRCLKX Q[3] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI6 D[4] DCTRCLK DCTRCLKX Q[4] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI7 D[5] DCTRCLK DCTRCLKX Q[5] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI8 D[6] DCTRCLK DCTRCLKX Q[6] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI9 D[7] DCTRCLK DCTRCLKX Q[7] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+STWL VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1_MD
XI10 D[8] DCTRCLK DCTRCLKX Q[8] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+VSS VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI11 D[9] DCTRCLK DCTRCLKX Q[9] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+VSS VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI12 D[10] DCTRCLK DCTRCLKX Q[10] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+VSS VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI13 D[11] DCTRCLK DCTRCLKX Q[11] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+VSS VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI14 D[12] DCTRCLK DCTRCLKX Q[12] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+VSS VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI15 D[13] DCTRCLK DCTRCLKX Q[13] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+VSS VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI16 D[14] DCTRCLK DCTRCLKX Q[14] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+VSS VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI17 D[15] DCTRCLK DCTRCLKX Q[15] RWLL[1] RWLL[0] RWLU[1] RWLU[0] SACK1 SACK4
+VSS VDD VSS WE WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256]
+WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_Y16_X512_D1
XI18 RWLU[0] RWLU[1] VDD VSS WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_PCAP_EDGE256_UP
XI19 RWLU[0] RWLU[1] VDD VSS WL[511] WL[510] WL[509] WL[508] WL[507] WL[506]
+WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496]
+WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486]
+WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476]
+WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466]
+WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456]
+WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446]
+WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436]
+WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426]
+WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416]
+WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406]
+WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396]
+WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386]
+WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376]
+WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366]
+WL[365] WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356]
+WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346]
+WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336]
+WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326]
+WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316]
+WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306]
+WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296]
+WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286]
+WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276]
+WL[275] WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266]
+WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256] S55NLLGSPH_X512Y16D32_PCAP_EDGE256_UP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_TIE_LOW_S
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_TIE_LOW_S PULL0 VSS VDD
MP18 VDD NET2 NET2 VDD P12LL W=2U L=0.06U M=1
MN18 PULL0 NET2 VSS VSS N12LL W=3U L=0.06U M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_TIE_HIGH_S
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_TIE_HIGH_S PULL1 VSS VDD
MP18 VDD NET2 PULL1 VDD P12LL W=4U L=0.06U M=1
MN18 NET2 NET2 VSS VSS N12LL W=2U L=0.06U M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_SOP_S
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_SOP_S DBL EMCLK S[1] S[0] VDD VSS
M0 9 8 VSS VSS N12LL L=6E-08 W=4E-07 $X=22095 $Y=1405 $D=0
M1 VSS 10 9 VSS N12LL L=6E-08 W=4E-07 $X=22385 $Y=1405 $D=0
M2 11 10 VSS VSS N12LL L=6E-08 W=4E-07 $X=22685 $Y=1405 $D=0
M3 43 10 12 VSS N12LL L=6E-08 W=4E-07 $X=23600 $Y=1490 $D=0
M4 VSS 8 43 VSS N12LL L=6E-08 W=4E-07 $X=23890 $Y=1490 $D=0
M5 S[1] VSS VSS VSS N12LL L=6E-08 W=2E-07 $X=24510 $Y=1630 $D=0
M6 VSS S[1] 10 VSS N12LL L=6E-08 W=4E-07 $X=25095 $Y=1420 $D=0
M7 8 S[0] VSS VSS N12LL L=6E-08 W=4E-07 $X=25385 $Y=1420 $D=0
M8 VSS VSS S[0] VSS N12LL L=6E-08 W=2E-07 $X=25980 $Y=1610 $D=0
M9 4 EMCLK DBL VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=16655 $Y=1555 $D=73
M10 4 EMCLK DBL VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=16655 $Y=1840 $D=73
M11 4 EMCLK DBL VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=16655 $Y=2345 $D=73
M12 4 EMCLK DBL VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=16655 $Y=2630 $D=73
M13 DBL EMCLK 5 VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=17760 $Y=1555 $D=73
M14 DBL EMCLK 5 VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=17760 $Y=1840 $D=73
M15 DBL EMCLK 5 VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=17760 $Y=2345 $D=73
M16 DBL EMCLK 5 VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=17760 $Y=2630 $D=73
M17 6 EMCLK DBL VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=18135 $Y=1555 $D=73
M18 6 EMCLK DBL VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=18135 $Y=1840 $D=73
M19 6 EMCLK DBL VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=18135 $Y=2345 $D=73
M20 6 EMCLK DBL VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=18135 $Y=2630 $D=73
M21 DBL EMCLK 7 VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=19240 $Y=1555 $D=73
M22 DBL EMCLK 7 VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=19240 $Y=1840 $D=73
M23 DBL EMCLK 7 VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=19240 $Y=2345 $D=73
M24 DBL EMCLK 7 VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=19240 $Y=2630 $D=73
M25 7 EMCLK DBL VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=19615 $Y=1555 $D=73
M26 7 EMCLK DBL VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=19615 $Y=1840 $D=73
M27 7 EMCLK DBL VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=19615 $Y=2345 $D=73
M28 7 EMCLK DBL VSS STNPGHVT W=8.5E-08 L=7.5E-08 $X=19615 $Y=2630 $D=73
M29 VSS VDD 4 VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=17020 $Y=1505 $D=72
M30 VSS VDD 4 VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=17020 $Y=1840 $D=72
M31 VSS VDD 4 VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=17020 $Y=2295 $D=72
M32 VSS VDD 4 VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=17020 $Y=2630 $D=72
M33 5 12 VSS VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=17405 $Y=1505 $D=72
M34 5 12 VSS VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=17405 $Y=1840 $D=72
M35 5 12 VSS VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=17405 $Y=2295 $D=72
M36 5 12 VSS VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=17405 $Y=2630 $D=72
M37 VSS 11 6 VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=18500 $Y=1505 $D=72
M38 VSS 11 6 VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=18500 $Y=1840 $D=72
M39 VSS 11 6 VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=18500 $Y=2295 $D=72
M40 VSS 11 6 VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=18500 $Y=2630 $D=72
M41 7 9 VSS VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=18885 $Y=1505 $D=72
M42 7 9 VSS VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=18885 $Y=1840 $D=72
M43 7 9 VSS VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=18885 $Y=2295 $D=72
M44 7 9 VSS VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=18885 $Y=2630 $D=72
M45 VSS 9 7 VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=19980 $Y=1505 $D=72
M46 VSS 9 7 VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=19980 $Y=1840 $D=72
M47 VSS 9 7 VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=19980 $Y=2295 $D=72
M48 VSS 9 7 VSS STNPDHVT W=1.35E-07 L=6.5E-08 $X=19980 $Y=2630 $D=72
M49 44 8 9 VDD P12LL L=6E-08 W=4E-07 $X=22165 $Y=2680 $D=2
M50 VDD 10 44 VDD P12LL L=6E-08 W=4E-07 $X=22385 $Y=2680 $D=2
M51 11 10 VDD VDD P12LL L=6E-08 W=4E-07 $X=22685 $Y=2680 $D=2
M52 12 10 VDD VDD P12LL L=6E-08 W=4E-07 $X=23600 $Y=2675 $D=2
M53 VDD 8 12 VDD P12LL L=6E-08 W=4E-07 $X=23890 $Y=2675 $D=2
M54 S[1] VDD VDD VDD P12LL L=6E-08 W=2E-07 $X=24510 $Y=2530 $D=2
M55 VDD S[1] 10 VDD P12LL L=6E-08 W=4E-07 $X=25095 $Y=2530 $D=2
M56 8 S[0] VDD VDD P12LL L=6E-08 W=4E-07 $X=25385 $Y=2530 $D=2
M57 VDD VDD S[0] VDD P12LL L=6E-08 W=2E-07 $X=25980 $Y=2530 $D=2
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_LOGIC_LEAFCELL_COMMON
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_LOGIC_LEAFCELL_COMMON RWLL RDE ACTRCLK ACTRCLKX ZAX PXA[3] PXA[2] PXA[1] PXA[0] XA[4]
+XA[3] XA[2] XA[1] XA[0] ZA FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3]
+FCKX[2] FCKX[1] FCKX[0] S[1] S[0] WEN WE CEN CLK FB
+YX[7] YX[6] YX[5] YX[4] YX[3] YX[2] YX[1] YX[0] YA[2] YA[1]
+YA[0] EMCLK RWLR SACK1 SACK4 DCTRCLK DCTRCLKX VDD VSS
M0 123 XA[3] VSS VSS N12LL L=6E-08 W=4E-07 $X=640 $Y=3130 $D=0
M1 VSS RDE 123 VSS N12LL L=6E-08 W=4E-07 $X=910 $Y=3130 $D=0
M2 124 123 VSS VSS N12LL L=3E-07 W=4E-07 $X=1220 $Y=3130 $D=0
M3 128 ZAX VSS VSS N12LL L=6E-07 W=1.2E-07 $X=1450 $Y=4420 $D=0
M4 VSS 124 125 VSS N12LL L=6E-08 W=4E-07 $X=2080 $Y=3130 $D=0
M5 127 125 VSS VSS N12LL L=6E-08 W=1E-06 $X=2400 $Y=3130 $D=0
M6 127 ACTRCLKX 128 VSS N12LL L=6E-08 W=1.245E-06 $X=3115 $Y=3130 $D=0
M7 128 ACTRCLKX 127 VSS N12LL L=6E-08 W=1.245E-06 $X=3385 $Y=3130 $D=0
M8 RWLL 131 VSS VSS N12LL L=6E-08 W=1E-06 $X=3940 $Y=33805 $D=0
M9 VSS 131 RWLL VSS N12LL L=6E-08 W=1E-06 $X=3940 $Y=34075 $D=0
M10 ZAX 128 VSS VSS N12LL L=6E-08 W=1.25E-06 $X=3995 $Y=3130 $D=0
M11 VSS 128 ZAX VSS N12LL L=6E-08 W=1.25E-06 $X=4265 $Y=3130 $D=0
M12 ZAX 128 VSS VSS N12LL L=6E-08 W=1.25E-06 $X=4535 $Y=3130 $D=0
M13 VSS 128 ZAX VSS N12LL L=6E-08 W=1.25E-06 $X=4805 $Y=3130 $D=0
M14 PXA[3] 132 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=5015 $Y=24970 $D=0
M15 142 134 VSS VSS N12LL L=6E-08 W=5E-07 $X=5095 $Y=11630 $D=0
M16 136 PXA[2] VSS VSS N12LL L=6E-07 W=1.2E-07 $X=5095 $Y=24185 $D=0
M17 133 128 VSS VSS N12LL L=6E-08 W=1E-06 $X=5115 $Y=3130 $D=0
M18 307 142 130 VSS N12LL L=6E-08 W=1.5E-06 $X=5130 $Y=13175 $D=0
M19 132 ACTRCLKX 130 VSS N12LL L=6E-08 W=2.5E-06 $X=5160 $Y=17420 $D=0
M20 VSS PXA[3] 132 VSS N12LL L=6E-07 W=1.2E-07 $X=5265 $Y=23500 $D=0
M21 VSS 132 PXA[3] VSS N12LL L=6E-08 W=1.5E-06 $X=5305 $Y=24970 $D=0
M22 VSS 140 307 VSS N12LL L=6E-08 W=1.5E-06 $X=5320 $Y=13175 $D=0
M23 VSS RDE 142 VSS N12LL L=6E-08 W=5E-07 $X=5385 $Y=11630 $D=0
M24 VSS XA[3] 134 VSS N12LL L=6E-08 W=4E-07 $X=5440 $Y=7445 $D=0
M25 131 209 58 VSS N12LL L=6E-08 W=1E-06 $X=5500 $Y=33805 $D=0
M26 308 140 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=5580 $Y=13175 $D=0
M27 PXA[2] 136 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=5595 $Y=24970 $D=0
M28 73 RDE VSS VSS N12LL L=6E-08 W=7E-07 $X=5675 $Y=11630 $D=0
M29 ZA 133 VSS VSS N12LL L=6E-08 W=1.25E-06 $X=5735 $Y=3130 $D=0
M30 135 ACTRCLKX 136 VSS N12LL L=6E-08 W=2.5E-06 $X=5740 $Y=17420 $D=0
M31 137 134 VSS VSS N12LL L=6E-08 W=4E-07 $X=5765 $Y=7445 $D=0
M32 135 73 308 VSS N12LL L=6E-08 W=1.5E-06 $X=5770 $Y=13175 $D=0
M33 VSS 136 PXA[2] VSS N12LL L=6E-08 W=1.5E-06 $X=5885 $Y=24970 $D=0
M34 VSS 137 73 VSS N12LL L=6E-08 W=7E-07 $X=5965 $Y=11630 $D=0
M35 VSS 133 ZA VSS N12LL L=6E-08 W=1.25E-06 $X=6005 $Y=3130 $D=0
M36 PXA[0] 138 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=6225 $Y=24970 $D=0
M37 ZA 133 VSS VSS N12LL L=6E-08 W=1.25E-06 $X=6275 $Y=3130 $D=0
M38 141 PXA[1] VSS VSS N12LL L=6E-07 W=1.2E-07 $X=6305 $Y=23500 $D=0
M39 309 73 139 VSS N12LL L=6E-08 W=1.5E-06 $X=6340 $Y=13175 $D=0
M40 138 ACTRCLKX 139 VSS N12LL L=6E-08 W=2.5E-06 $X=6370 $Y=17420 $D=0
M41 VSS PXA[0] 138 VSS N12LL L=6E-07 W=1.2E-07 $X=6475 $Y=24185 $D=0
M42 310 VDD VSS VSS N12LL L=3E-07 W=4E-07 $X=6480 $Y=7445 $D=0
M43 VSS 138 PXA[0] VSS N12LL L=6E-08 W=1.5E-06 $X=6515 $Y=24970 $D=0
M44 VSS 145 309 VSS N12LL L=6E-08 W=1.5E-06 $X=6530 $Y=13175 $D=0
M45 VSS 133 ZA VSS N12LL L=6E-08 W=1.25E-06 $X=6545 $Y=3130 $D=0
M46 311 145 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=6790 $Y=13175 $D=0
M47 PXA[1] 141 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=6805 $Y=24970 $D=0
M48 VSS 144 140 VSS N12LL L=6E-08 W=7E-07 $X=6820 $Y=11630 $D=0
M49 143 ACTRCLKX 141 VSS N12LL L=6E-08 W=2.5E-06 $X=6950 $Y=17420 $D=0
M50 143 142 311 VSS N12LL L=6E-08 W=1.5E-06 $X=6980 $Y=13175 $D=0
M51 144 XA[4] 310 VSS N12LL L=6E-08 W=4E-07 $X=7000 $Y=7445 $D=0
M52 VSS 141 PXA[1] VSS N12LL L=6E-08 W=1.5E-06 $X=7095 $Y=24970 $D=0
M53 145 140 VSS VSS N12LL L=6E-08 W=7E-07 $X=7110 $Y=11630 $D=0
M54 76 149 VSS VSS N12LL L=6E-08 W=4E-07 $X=8705 $Y=25095 $D=0
M55 FCKX[3] 76 58 VSS N12LL L=6E-08 W=1.25E-06 $X=8705 $Y=29015 $D=0
M56 161 188 VSS VSS N12LL L=6E-08 W=5E-07 $X=8865 $Y=15060 $D=0
M57 152 ACTRCLKX 149 VSS N12LL L=6E-08 W=5E-07 $X=8865 $Y=21055 $D=0
M58 VSS 76 149 VSS N12LL L=6E-07 W=1.2E-07 $X=8955 $Y=26265 $D=0
M59 VSS 149 76 VSS N12LL L=6E-08 W=4E-07 $X=8995 $Y=25095 $D=0
M60 58 76 FCKX[3] VSS N12LL L=6E-08 W=1.25E-06 $X=8995 $Y=29015 $D=0
M61 312 61 152 VSS N12LL L=6E-08 W=1E-06 $X=9095 $Y=19480 $D=0
M62 VSS 188 161 VSS N12LL L=6E-08 W=5E-07 $X=9135 $Y=15060 $D=0
M63 149 ACTRCLKX 152 VSS N12LL L=6E-08 W=5E-07 $X=9135 $Y=21055 $D=0
M64 76 149 VSS VSS N12LL L=6E-08 W=4E-07 $X=9285 $Y=25095 $D=0
M65 FCKX[3] 76 58 VSS N12LL L=6E-08 W=1.25E-06 $X=9285 $Y=29015 $D=0
M66 313 60 312 VSS N12LL L=6E-08 W=1E-06 $X=9335 $Y=19480 $D=0
M67 152 ACTRCLKX 149 VSS N12LL L=6E-08 W=5E-07 $X=9415 $Y=21055 $D=0
M68 188 155 VSS VSS N12LL L=6E-08 W=5E-07 $X=9425 $Y=15060 $D=0
M69 VSS 161 313 VSS N12LL L=6E-08 W=1E-06 $X=9575 $Y=19480 $D=0
M70 VSS 149 76 VSS N12LL L=6E-08 W=4E-07 $X=9575 $Y=25095 $D=0
M71 58 76 FCKX[3] VSS N12LL L=6E-08 W=1.25E-06 $X=9575 $Y=29015 $D=0
M72 VSS 155 188 VSS N12LL L=6E-08 W=5E-07 $X=9715 $Y=15060 $D=0
M73 314 161 VSS VSS N12LL L=6E-08 W=1E-06 $X=9865 $Y=19480 $D=0
M74 80 156 VSS VSS N12LL L=6E-08 W=4E-07 $X=9865 $Y=25095 $D=0
M75 FCKX[2] 80 58 VSS N12LL L=6E-08 W=1.25E-06 $X=9865 $Y=29015 $D=0
M76 156 80 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=9945 $Y=26265 $D=0
M77 156 ACTRCLKX 78 VSS N12LL L=6E-08 W=5E-07 $X=10025 $Y=21055 $D=0
M78 315 60 314 VSS N12LL L=6E-08 W=1E-06 $X=10105 $Y=19480 $D=0
M79 VSS 156 80 VSS N12LL L=6E-08 W=4E-07 $X=10155 $Y=25095 $D=0
M80 58 80 FCKX[2] VSS N12LL L=6E-08 W=1.25E-06 $X=10155 $Y=29015 $D=0
M81 78 ACTRCLKX 156 VSS N12LL L=6E-08 W=5E-07 $X=10305 $Y=21055 $D=0
M82 316 XA[2] 155 VSS N12LL L=6E-08 W=4E-07 $X=10345 $Y=15140 $D=0
M83 78 59 315 VSS N12LL L=6E-08 W=1E-06 $X=10345 $Y=19480 $D=0
M84 80 156 VSS VSS N12LL L=6E-08 W=4E-07 $X=10445 $Y=25095 $D=0
M85 FCKX[2] 80 58 VSS N12LL L=6E-08 W=1.25E-06 $X=10445 $Y=29015 $D=0
M86 VSS VDD 316 VSS N12LL L=3E-07 W=4E-07 $X=10575 $Y=15140 $D=0
M87 156 ACTRCLKX 78 VSS N12LL L=6E-08 W=5E-07 $X=10575 $Y=21055 $D=0
M88 VSS 156 80 VSS N12LL L=6E-08 W=4E-07 $X=10735 $Y=25095 $D=0
M89 58 80 FCKX[2] VSS N12LL L=6E-08 W=1.25E-06 $X=10735 $Y=29015 $D=0
M90 185 198 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=10825 $Y=33505 $D=0
M91 82 160 VSS VSS N12LL L=6E-08 W=4E-07 $X=11025 $Y=25095 $D=0
M92 FCKX[0] 82 58 VSS N12LL L=6E-08 W=1.25E-06 $X=11025 $Y=29015 $D=0
M93 84 ACTRCLKX 160 VSS N12LL L=6E-08 W=5E-07 $X=11185 $Y=21055 $D=0
M94 VSS 82 160 VSS N12LL L=6E-07 W=1.2E-07 $X=11275 $Y=26265 $D=0
M95 VSS 160 82 VSS N12LL L=6E-08 W=4E-07 $X=11315 $Y=25095 $D=0
M96 58 82 FCKX[0] VSS N12LL L=6E-08 W=1.25E-06 $X=11315 $Y=29015 $D=0
M97 318 59 84 VSS N12LL L=6E-08 W=1E-06 $X=11415 $Y=19480 $D=0
M98 160 ACTRCLKX 84 VSS N12LL L=6E-08 W=5E-07 $X=11455 $Y=21055 $D=0
M99 82 160 VSS VSS N12LL L=6E-08 W=4E-07 $X=11605 $Y=25095 $D=0
M100 FCKX[0] 82 58 VSS N12LL L=6E-08 W=1.25E-06 $X=11605 $Y=29015 $D=0
M101 319 194 318 VSS N12LL L=6E-08 W=1E-06 $X=11655 $Y=19480 $D=0
M102 320 162 83 VSS N12LL L=6E-08 W=4E-07 $X=11690 $Y=12335 $D=0
M103 84 ACTRCLKX 160 VSS N12LL L=6E-08 W=5E-07 $X=11735 $Y=21055 $D=0
M104 VSS S[0] 162 VSS N12LL L=6E-08 W=4E-07 $X=11790 $Y=10790 $D=0
M105 VSS 161 319 VSS N12LL L=6E-08 W=1E-06 $X=11895 $Y=19480 $D=0
M106 VSS 160 82 VSS N12LL L=6E-08 W=4E-07 $X=11895 $Y=25095 $D=0
M107 58 82 FCKX[0] VSS N12LL L=6E-08 W=1.25E-06 $X=11895 $Y=29015 $D=0
M108 VSS 88 320 VSS N12LL L=6E-08 W=4E-07 $X=11960 $Y=12335 $D=0
M109 164 WEN VSS VSS N12LL L=6E-08 W=4E-07 $X=11990 $Y=1520 $D=0
M110 173 162 VSS VSS N12LL L=6E-08 W=4E-07 $X=12060 $Y=10790 $D=0
M111 85 163 VSS VSS N12LL L=6E-08 W=1E-06 $X=12145 $Y=4990 $D=0
M112 321 161 VSS VSS N12LL L=6E-08 W=1E-06 $X=12185 $Y=19480 $D=0
M113 86 165 VSS VSS N12LL L=6E-08 W=4E-07 $X=12185 $Y=25095 $D=0
M114 FCKX[1] 86 58 VSS N12LL L=6E-08 W=1.25E-06 $X=12185 $Y=29015 $D=0
M115 208 83 VSS VSS N12LL L=6E-08 W=4E-07 $X=12230 $Y=12335 $D=0
M116 185 ACTRCLKX 176 VSS N12LL L=6E-08 W=1E-06 $X=12255 $Y=33930 $D=0
M117 165 86 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=12265 $Y=26265 $D=0
M118 165 ACTRCLKX 166 VSS N12LL L=6E-08 W=5E-07 $X=12345 $Y=21055 $D=0
M119 323 VDD VSS VSS N12LL L=3E-07 W=4E-07 $X=12405 $Y=15140 $D=0
M120 322 194 321 VSS N12LL L=6E-08 W=1E-06 $X=12425 $Y=19480 $D=0
M121 VSS 165 86 VSS N12LL L=6E-08 W=4E-07 $X=12475 $Y=25095 $D=0
M122 58 86 FCKX[1] VSS N12LL L=6E-08 W=1.25E-06 $X=12475 $Y=29015 $D=0
M123 166 ACTRCLKX 165 VSS N12LL L=6E-08 W=5E-07 $X=12625 $Y=21055 $D=0
M124 324 85 168 VSS N12LL L=6E-08 W=3E-06 $X=12655 $Y=2990 $D=0
M125 166 61 322 VSS N12LL L=6E-08 W=1E-06 $X=12665 $Y=19480 $D=0
M126 VSS 164 167 VSS N12LL L=3E-07 W=4E-07 $X=12695 $Y=1520 $D=0
M127 VSS 185 198 VSS N12LL L=6E-08 W=4E-07 $X=12695 $Y=34560 $D=0
M128 209 198 VSS VSS N12LL L=6E-08 W=4E-07 $X=12695 $Y=34830 $D=0
M129 86 165 VSS VSS N12LL L=6E-08 W=4E-07 $X=12765 $Y=25095 $D=0
M130 FCKX[1] 86 58 VSS N12LL L=6E-08 W=1.25E-06 $X=12765 $Y=29015 $D=0
M131 VSS RDE 182 VSS N12LL L=6E-08 W=4E-07 $X=12855 $Y=33350 $D=0
M132 176 182 VSS VSS N12LL L=6E-08 W=4E-07 $X=12855 $Y=33620 $D=0
M133 VSS 49 324 VSS N12LL L=6E-08 W=3E-06 $X=12875 $Y=2990 $D=0
M134 169 XA[0] 323 VSS N12LL L=6E-08 W=4E-07 $X=12875 $Y=15140 $D=0
M135 165 ACTRCLKX 166 VSS N12LL L=6E-08 W=5E-07 $X=12895 $Y=21055 $D=0
M136 325 173 87 VSS N12LL L=6E-08 W=4E-07 $X=12920 $Y=12290 $D=0
M137 VSS 165 86 VSS N12LL L=6E-08 W=4E-07 $X=13055 $Y=25095 $D=0
M138 58 86 FCKX[1] VSS N12LL L=6E-08 W=1.25E-06 $X=13055 $Y=29015 $D=0
M139 WE 168 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=13125 $Y=3490 $D=0
M140 VSS 85 163 VSS N12LL L=6E-07 W=1.2E-07 $X=13165 $Y=2465 $D=0
M141 VSS 174 325 VSS N12LL L=6E-08 W=4E-07 $X=13260 $Y=12290 $D=0
M142 171 167 VSS VSS N12LL L=2E-07 W=4E-07 $X=13325 $Y=1520 $D=0
M143 89 170 VSS VSS N12LL L=6E-08 W=4E-07 $X=13345 $Y=25095 $D=0
M144 FCKX[7] 89 58 VSS N12LL L=6E-08 W=1.25E-06 $X=13345 $Y=29015 $D=0
M145 VSS 168 WE VSS N12LL L=6E-08 W=2.5E-06 $X=13375 $Y=3490 $D=0
M146 VSS S[1] 174 VSS N12LL L=6E-08 W=4E-07 $X=13405 $Y=10910 $D=0
M147 61 169 VSS VSS N12LL L=6E-08 W=5E-07 $X=13505 $Y=15060 $D=0
M148 90 ACTRCLKX 170 VSS N12LL L=6E-08 W=5E-07 $X=13505 $Y=21055 $D=0
M149 172 87 VSS VSS N12LL L=6E-08 W=4E-07 $X=13530 $Y=12290 $D=0
M150 VSS 89 170 VSS N12LL L=6E-07 W=1.2E-07 $X=13595 $Y=26265 $D=0
M151 VSS 170 89 VSS N12LL L=6E-08 W=4E-07 $X=13635 $Y=25095 $D=0
M152 58 89 FCKX[7] VSS N12LL L=6E-08 W=1.25E-06 $X=13635 $Y=29015 $D=0
M153 88 174 VSS VSS N12LL L=6E-08 W=4E-07 $X=13665 $Y=10910 $D=0
M154 326 61 90 VSS N12LL L=6E-08 W=1E-06 $X=13735 $Y=19480 $D=0
M155 170 ACTRCLKX 90 VSS N12LL L=6E-08 W=5E-07 $X=13775 $Y=21055 $D=0
M156 VSS 169 61 VSS N12LL L=6E-08 W=5E-07 $X=13795 $Y=15060 $D=0
M157 89 170 VSS VSS N12LL L=6E-08 W=4E-07 $X=13925 $Y=25095 $D=0
M158 FCKX[7] 89 58 VSS N12LL L=6E-08 W=1.25E-06 $X=13925 $Y=29015 $D=0
M159 327 60 326 VSS N12LL L=6E-08 W=1E-06 $X=13975 $Y=19480 $D=0
M160 90 ACTRCLKX 170 VSS N12LL L=6E-08 W=5E-07 $X=14055 $Y=21055 $D=0
M161 59 61 VSS VSS N12LL L=6E-08 W=5E-07 $X=14085 $Y=15060 $D=0
M162 175 171 VSS VSS N12LL L=6E-08 W=1E-06 $X=14105 $Y=1585 $D=0
M163 328 162 181 VSS N12LL L=6E-08 W=4E-07 $X=14130 $Y=12290 $D=0
M164 VSS 188 327 VSS N12LL L=6E-08 W=1E-06 $X=14215 $Y=19480 $D=0
M165 VSS 170 89 VSS N12LL L=6E-08 W=4E-07 $X=14215 $Y=25095 $D=0
M166 58 89 FCKX[7] VSS N12LL L=6E-08 W=1.25E-06 $X=14215 $Y=29015 $D=0
M167 329 173 183 VSS N12LL L=6E-08 W=4E-07 $X=14260 $Y=10855 $D=0
M168 VSS 61 59 VSS N12LL L=6E-08 W=5E-07 $X=14355 $Y=15060 $D=0
M169 163 ACTRCLKX 175 VSS N12LL L=6E-08 W=1E-06 $X=14375 $Y=1585 $D=0
M170 VSS 174 328 VSS N12LL L=6E-08 W=4E-07 $X=14400 $Y=12290 $D=0
M171 VSS 177 196 VSS N12LL L=6E-08 W=2.5E-06 $X=14415 $Y=3490 $D=0
M172 330 188 VSS VSS N12LL L=6E-08 W=1E-06 $X=14505 $Y=19480 $D=0
M173 92 180 VSS VSS N12LL L=6E-08 W=4E-07 $X=14505 $Y=25095 $D=0
M174 FCKX[6] 92 58 VSS N12LL L=6E-08 W=1.25E-06 $X=14505 $Y=29015 $D=0
M175 VSS 88 329 VSS N12LL L=6E-08 W=4E-07 $X=14530 $Y=10855 $D=0
M176 180 92 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=14585 $Y=26265 $D=0
M177 180 ACTRCLKX 91 VSS N12LL L=6E-08 W=5E-07 $X=14665 $Y=21055 $D=0
M178 178 181 VSS VSS N12LL L=6E-08 W=4E-07 $X=14670 $Y=12290 $D=0
M179 177 FB VSS VSS N12LL L=6E-08 W=8E-07 $X=14745 $Y=5190 $D=0
M180 331 60 330 VSS N12LL L=6E-08 W=1E-06 $X=14745 $Y=19480 $D=0
M181 VSS 180 92 VSS N12LL L=6E-08 W=4E-07 $X=14795 $Y=25095 $D=0
M182 58 92 FCKX[6] VSS N12LL L=6E-08 W=1.25E-06 $X=14795 $Y=29015 $D=0
M183 184 183 VSS VSS N12LL L=6E-08 W=4E-07 $X=14800 $Y=10855 $D=0
M184 91 ACTRCLKX 180 VSS N12LL L=6E-08 W=5E-07 $X=14945 $Y=21055 $D=0
M185 VSS CLK 179 VSS N12LL L=6E-08 W=4E-07 $X=14955 $Y=1500 $D=0
M186 91 59 331 VSS N12LL L=6E-08 W=1E-06 $X=14985 $Y=19480 $D=0
M187 92 180 VSS VSS N12LL L=6E-08 W=4E-07 $X=15085 $Y=25095 $D=0
M188 FCKX[6] 92 58 VSS N12LL L=6E-08 W=1.25E-06 $X=15085 $Y=29015 $D=0
M189 180 ACTRCLKX 91 VSS N12LL L=6E-08 W=5E-07 $X=15215 $Y=21055 $D=0
M190 332 179 VSS VSS N12LL L=6E-08 W=1E-06 $X=15305 $Y=1500 $D=0
M191 VSS CLK 204 VSS N12LL L=6E-08 W=2.5E-06 $X=15330 $Y=3490 $D=0
M192 VSS 180 92 VSS N12LL L=6E-08 W=4E-07 $X=15375 $Y=25095 $D=0
M193 58 92 FCKX[6] VSS N12LL L=6E-08 W=1.25E-06 $X=15375 $Y=29015 $D=0
M194 190 CEN 332 VSS N12LL L=6E-08 W=1E-06 $X=15545 $Y=1500 $D=0
M195 333 VDD VSS VSS N12LL L=3E-07 W=4E-07 $X=15585 $Y=15140 $D=0
M196 204 CLK VSS VSS N12LL L=6E-08 W=2.5E-06 $X=15600 $Y=3490 $D=0
M197 93 186 VSS VSS N12LL L=6E-08 W=4E-07 $X=15665 $Y=25095 $D=0
M198 FCKX[4] 93 58 VSS N12LL L=6E-08 W=1.25E-06 $X=15665 $Y=29015 $D=0
M199 94 ACTRCLKX 186 VSS N12LL L=6E-08 W=5E-07 $X=15825 $Y=21055 $D=0
M200 EMCLK 178 187 VSS N12LL L=6E-08 W=1.25E-06 $X=15860 $Y=12210 $D=0
M201 VSS CLK 204 VSS N12LL L=6E-08 W=2.5E-06 $X=15870 $Y=3490 $D=0
M202 VSS 192 190 VSS N12LL L=6E-07 W=1.2E-07 $X=15905 $Y=1635 $D=0
M203 VSS 93 186 VSS N12LL L=6E-07 W=1.2E-07 $X=15915 $Y=26265 $D=0
M204 VSS 186 93 VSS N12LL L=6E-08 W=4E-07 $X=15955 $Y=25095 $D=0
M205 58 93 FCKX[4] VSS N12LL L=6E-08 W=1.25E-06 $X=15955 $Y=29015 $D=0
M206 189 XA[1] 333 VSS N12LL L=6E-08 W=4E-07 $X=16055 $Y=15140 $D=0
M207 334 59 94 VSS N12LL L=6E-08 W=1E-06 $X=16055 $Y=19480 $D=0
M208 186 ACTRCLKX 94 VSS N12LL L=6E-08 W=5E-07 $X=16095 $Y=21055 $D=0
M209 187 178 EMCLK VSS N12LL L=6E-08 W=1.25E-06 $X=16130 $Y=12210 $D=0
M210 204 CLK VSS VSS N12LL L=6E-08 W=2.5E-06 $X=16140 $Y=3490 $D=0
M211 93 186 VSS VSS N12LL L=6E-08 W=4E-07 $X=16245 $Y=25095 $D=0
M212 FCKX[4] 93 58 VSS N12LL L=6E-08 W=1.25E-06 $X=16245 $Y=29015 $D=0
M213 335 194 334 VSS N12LL L=6E-08 W=1E-06 $X=16295 $Y=19480 $D=0
M214 94 ACTRCLKX 186 VSS N12LL L=6E-08 W=5E-07 $X=16375 $Y=21055 $D=0
M215 VSS CLK 204 VSS N12LL L=6E-08 W=2.5E-06 $X=16410 $Y=3490 $D=0
M216 VSS 191 187 VSS N12LL L=6E-08 W=7E-07 $X=16460 $Y=12210 $D=0
M217 VSS 188 335 VSS N12LL L=6E-08 W=1E-06 $X=16535 $Y=19480 $D=0
M218 VSS 186 93 VSS N12LL L=6E-08 W=4E-07 $X=16535 $Y=25095 $D=0
M219 58 93 FCKX[4] VSS N12LL L=6E-08 W=1.25E-06 $X=16535 $Y=29015 $D=0
M220 204 CLK VSS VSS N12LL L=6E-08 W=2.5E-06 $X=16680 $Y=3490 $D=0
M221 60 189 VSS VSS N12LL L=6E-08 W=5E-07 $X=16685 $Y=15060 $D=0
M222 336 188 VSS VSS N12LL L=6E-08 W=1E-06 $X=16825 $Y=19480 $D=0
M223 96 193 VSS VSS N12LL L=6E-08 W=4E-07 $X=16825 $Y=25095 $D=0
M224 FCKX[5] 96 58 VSS N12LL L=6E-08 W=1.25E-06 $X=16825 $Y=29015 $D=0
M225 192 190 VSS VSS N12LL L=6E-08 W=4E-07 $X=16835 $Y=1635 $D=0
M226 193 96 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=16905 $Y=26265 $D=0
M227 VSS CLK 204 VSS N12LL L=6E-08 W=2.5E-06 $X=16950 $Y=3490 $D=0
M228 VSS 189 60 VSS N12LL L=6E-08 W=5E-07 $X=16975 $Y=15060 $D=0
M229 193 ACTRCLKX 195 VSS N12LL L=6E-08 W=5E-07 $X=16985 $Y=21055 $D=0
M230 337 194 336 VSS N12LL L=6E-08 W=1E-06 $X=17065 $Y=19480 $D=0
M231 VSS 193 96 VSS N12LL L=6E-08 W=4E-07 $X=17115 $Y=25095 $D=0
M232 58 96 FCKX[5] VSS N12LL L=6E-08 W=1.25E-06 $X=17115 $Y=29015 $D=0
M233 204 CLK VSS VSS N12LL L=6E-08 W=2.5E-06 $X=17220 $Y=3490 $D=0
M234 194 60 VSS VSS N12LL L=6E-08 W=5E-07 $X=17265 $Y=15060 $D=0
M235 195 ACTRCLKX 193 VSS N12LL L=6E-08 W=5E-07 $X=17265 $Y=21055 $D=0
M236 195 61 337 VSS N12LL L=6E-08 W=1E-06 $X=17305 $Y=19480 $D=0
M237 VSS 203 191 VSS N12LL L=3E-07 W=7E-07 $X=17320 $Y=12050 $D=0
M238 96 193 VSS VSS N12LL L=6E-08 W=4E-07 $X=17405 $Y=25095 $D=0
M239 FCKX[5] 96 58 VSS N12LL L=6E-08 W=1.25E-06 $X=17405 $Y=29015 $D=0
M240 197 192 VSS VSS N12LL L=6E-08 W=5E-07 $X=17445 $Y=1610 $D=0
M241 103 202 204 VSS N12LL L=6E-08 W=2.5E-06 $X=17490 $Y=3490 $D=0
M242 VSS 60 194 VSS N12LL L=6E-08 W=5E-07 $X=17535 $Y=15060 $D=0
M243 193 ACTRCLKX 195 VSS N12LL L=6E-08 W=5E-07 $X=17535 $Y=21055 $D=0
M244 VSS 193 96 VSS N12LL L=6E-08 W=4E-07 $X=17695 $Y=25095 $D=0
M245 58 96 FCKX[5] VSS N12LL L=6E-08 W=1.25E-06 $X=17695 $Y=29015 $D=0
M246 VSS CLK 197 VSS N12LL L=6E-08 W=5E-07 $X=17715 $Y=1610 $D=0
M247 204 202 103 VSS N12LL L=6E-08 W=2.5E-06 $X=17760 $Y=3490 $D=0
M248 207 99 VSS VSS N12LL L=3E-07 W=7E-07 $X=17910 $Y=12050 $D=0
M249 200 197 VSS VSS N12LL L=6E-08 W=5E-07 $X=17985 $Y=1610 $D=0
M250 98 199 VSS VSS N12LL L=6E-08 W=4E-07 $X=17985 $Y=25095 $D=0
M251 YX[3] 98 58 VSS N12LL L=6E-08 W=1.25E-06 $X=17985 $Y=29015 $D=0
M252 103 202 204 VSS N12LL L=6E-08 W=2.5E-06 $X=18030 $Y=3490 $D=0
M253 211 226 VSS VSS N12LL L=6E-08 W=5E-07 $X=18145 $Y=15060 $D=0
M254 201 ACTRCLKX 199 VSS N12LL L=6E-08 W=5E-07 $X=18145 $Y=21055 $D=0
M255 VSS 98 199 VSS N12LL L=6E-07 W=1.2E-07 $X=18235 $Y=26265 $D=0
M256 VSS 199 98 VSS N12LL L=6E-08 W=4E-07 $X=18275 $Y=25095 $D=0
M257 58 98 YX[3] VSS N12LL L=6E-08 W=1.25E-06 $X=18275 $Y=29015 $D=0
M258 204 202 103 VSS N12LL L=6E-08 W=2.5E-06 $X=18300 $Y=3490 $D=0
M259 338 71 201 VSS N12LL L=6E-08 W=1E-06 $X=18375 $Y=19480 $D=0
M260 VSS 226 211 VSS N12LL L=6E-08 W=5E-07 $X=18415 $Y=15060 $D=0
M261 199 ACTRCLKX 201 VSS N12LL L=6E-08 W=5E-07 $X=18415 $Y=21055 $D=0
M262 98 199 VSS VSS N12LL L=6E-08 W=4E-07 $X=18565 $Y=25095 $D=0
M263 YX[3] 98 58 VSS N12LL L=6E-08 W=1.25E-06 $X=18565 $Y=29015 $D=0
M264 103 202 204 VSS N12LL L=6E-08 W=2.5E-06 $X=18570 $Y=3490 $D=0
M265 202 200 VSS VSS N12LL L=6E-08 W=5E-07 $X=18595 $Y=1610 $D=0
M266 339 68 338 VSS N12LL L=6E-08 W=1E-06 $X=18615 $Y=19480 $D=0
M267 201 ACTRCLKX 199 VSS N12LL L=6E-08 W=5E-07 $X=18695 $Y=21055 $D=0
M268 226 205 VSS VSS N12LL L=6E-08 W=5E-07 $X=18705 $Y=15060 $D=0
M269 204 202 103 VSS N12LL L=6E-08 W=2.5E-06 $X=18840 $Y=3490 $D=0
M270 VSS 211 339 VSS N12LL L=6E-08 W=1E-06 $X=18855 $Y=19480 $D=0
M271 VSS 199 98 VSS N12LL L=6E-08 W=4E-07 $X=18855 $Y=25095 $D=0
M272 58 98 YX[3] VSS N12LL L=6E-08 W=1.25E-06 $X=18855 $Y=29015 $D=0
M273 VSS 200 202 VSS N12LL L=6E-08 W=5E-07 $X=18865 $Y=1610 $D=0
M274 VSS 205 226 VSS N12LL L=6E-08 W=5E-07 $X=18995 $Y=15060 $D=0
M275 103 202 204 VSS N12LL L=6E-08 W=2.5E-06 $X=19110 $Y=3490 $D=0
M276 EMCLK 172 203 VSS N12LL L=6E-08 W=1.25E-06 $X=19115 $Y=12050 $D=0
M277 202 200 VSS VSS N12LL L=6E-08 W=5E-07 $X=19135 $Y=1610 $D=0
M278 340 211 VSS VSS N12LL L=6E-08 W=1E-06 $X=19145 $Y=19480 $D=0
M279 101 206 VSS VSS N12LL L=6E-08 W=4E-07 $X=19145 $Y=25095 $D=0
M280 YX[2] 101 58 VSS N12LL L=6E-08 W=1.25E-06 $X=19145 $Y=29015 $D=0
M281 206 101 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=19225 $Y=26265 $D=0
M282 206 ACTRCLKX 102 VSS N12LL L=6E-08 W=5E-07 $X=19305 $Y=21055 $D=0
M283 203 172 EMCLK VSS N12LL L=6E-08 W=1.25E-06 $X=19365 $Y=12050 $D=0
M284 204 202 103 VSS N12LL L=6E-08 W=2.5E-06 $X=19380 $Y=3490 $D=0
M285 341 68 340 VSS N12LL L=6E-08 W=1E-06 $X=19385 $Y=19480 $D=0
M286 VSS 206 101 VSS N12LL L=6E-08 W=4E-07 $X=19435 $Y=25095 $D=0
M287 58 101 YX[2] VSS N12LL L=6E-08 W=1.25E-06 $X=19435 $Y=29015 $D=0
M288 102 ACTRCLKX 206 VSS N12LL L=6E-08 W=5E-07 $X=19585 $Y=21055 $D=0
M289 342 YA[2] 205 VSS N12LL L=6E-08 W=4E-07 $X=19625 $Y=15140 $D=0
M290 102 67 341 VSS N12LL L=6E-08 W=1E-06 $X=19625 $Y=19480 $D=0
M291 VSS 207 203 VSS N12LL L=6E-08 W=7E-07 $X=19710 $Y=12050 $D=0
M292 101 206 VSS VSS N12LL L=6E-08 W=4E-07 $X=19725 $Y=25095 $D=0
M293 YX[2] 101 58 VSS N12LL L=6E-08 W=1.25E-06 $X=19725 $Y=29015 $D=0
M294 VSS VDD 342 VSS N12LL L=3E-07 W=4E-07 $X=19855 $Y=15140 $D=0
M295 206 ACTRCLKX 102 VSS N12LL L=6E-08 W=5E-07 $X=19855 $Y=21055 $D=0
M296 49 103 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=19975 $Y=3590 $D=0
M297 99 212 VSS VSS N12LL L=6E-08 W=7E-07 $X=19980 $Y=12050 $D=0
M298 VSS 206 101 VSS N12LL L=6E-08 W=4E-07 $X=20015 $Y=25095 $D=0
M299 58 101 YX[2] VSS N12LL L=6E-08 W=1.25E-06 $X=20015 $Y=29015 $D=0
M300 VSS 49 103 VSS N12LL L=1E-06 W=1.2E-07 $X=20105 $Y=2765 $D=0
M301 VSS 213 220 VSS N12LL L=2E-07 W=4E-07 $X=20145 $Y=1805 $D=0
M302 VSS 103 49 VSS N12LL L=6E-08 W=2.5E-06 $X=20245 $Y=3590 $D=0
M303 105 210 VSS VSS N12LL L=6E-08 W=4E-07 $X=20305 $Y=25095 $D=0
M304 YX[0] 105 58 VSS N12LL L=6E-08 W=1.25E-06 $X=20305 $Y=29015 $D=0
M305 EMCLK 208 99 VSS N12LL L=6E-08 W=1.25E-06 $X=20320 $Y=12050 $D=0
M306 104 ACTRCLKX 210 VSS N12LL L=6E-08 W=5E-07 $X=20465 $Y=21055 $D=0
M307 49 103 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=20515 $Y=3590 $D=0
M308 VSS 105 210 VSS N12LL L=6E-07 W=1.2E-07 $X=20555 $Y=26265 $D=0
M309 99 208 EMCLK VSS N12LL L=6E-08 W=1.25E-06 $X=20570 $Y=12050 $D=0
M310 VSS 210 105 VSS N12LL L=6E-08 W=4E-07 $X=20595 $Y=25095 $D=0
M311 58 105 YX[0] VSS N12LL L=6E-08 W=1.25E-06 $X=20595 $Y=29015 $D=0
M312 213 VSS VSS VSS N12LL L=2E-07 W=4E-07 $X=20615 $Y=1805 $D=0
M313 343 67 104 VSS N12LL L=6E-08 W=1E-06 $X=20695 $Y=19480 $D=0
M314 210 ACTRCLKX 104 VSS N12LL L=6E-08 W=5E-07 $X=20735 $Y=21055 $D=0
M315 215 209 58 VSS N12LL L=6E-08 W=1E-06 $X=20750 $Y=33805 $D=0
M316 VSS 103 49 VSS N12LL L=6E-08 W=2.5E-06 $X=20785 $Y=3590 $D=0
M317 105 210 VSS VSS N12LL L=6E-08 W=4E-07 $X=20885 $Y=25095 $D=0
M318 YX[0] 105 58 VSS N12LL L=6E-08 W=1.25E-06 $X=20885 $Y=29015 $D=0
M319 344 230 343 VSS N12LL L=6E-08 W=1E-06 $X=20935 $Y=19480 $D=0
M320 104 ACTRCLKX 210 VSS N12LL L=6E-08 W=5E-07 $X=21015 $Y=21055 $D=0
M321 58 49 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=21075 $Y=3590 $D=0
M322 VSS 49 213 VSS N12LL L=2E-07 W=4E-07 $X=21105 $Y=1805 $D=0
M323 VSS 211 344 VSS N12LL L=6E-08 W=1E-06 $X=21175 $Y=19480 $D=0
M324 VSS 210 105 VSS N12LL L=6E-08 W=4E-07 $X=21175 $Y=25095 $D=0
M325 58 105 YX[0] VSS N12LL L=6E-08 W=1.25E-06 $X=21175 $Y=29015 $D=0
M326 VSS 218 212 VSS N12LL L=3E-07 W=7E-07 $X=21190 $Y=12050 $D=0
M327 VSS 49 58 VSS N12LL L=6E-08 W=2.5E-06 $X=21345 $Y=3590 $D=0
M328 345 211 VSS VSS N12LL L=6E-08 W=1E-06 $X=21465 $Y=19480 $D=0
M329 106 214 VSS VSS N12LL L=6E-08 W=4E-07 $X=21465 $Y=25095 $D=0
M330 YX[1] 106 58 VSS N12LL L=6E-08 W=1.25E-06 $X=21465 $Y=29015 $D=0
M331 214 106 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=21545 $Y=26265 $D=0
M332 58 49 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=21615 $Y=3590 $D=0
M333 214 ACTRCLKX 216 VSS N12LL L=6E-08 W=5E-07 $X=21625 $Y=21055 $D=0
M334 347 VDD VSS VSS N12LL L=3E-07 W=4E-07 $X=21685 $Y=15140 $D=0
M335 346 230 345 VSS N12LL L=6E-08 W=1E-06 $X=21705 $Y=19480 $D=0
M336 VSS 214 106 VSS N12LL L=6E-08 W=4E-07 $X=21755 $Y=25095 $D=0
M337 58 106 YX[1] VSS N12LL L=6E-08 W=1.25E-06 $X=21755 $Y=29015 $D=0
M338 VSS 49 58 VSS N12LL L=6E-08 W=2.5E-06 $X=21885 $Y=3590 $D=0
M339 VSS 49 217 VSS N12LL L=2E-07 W=4E-07 $X=21895 $Y=1805 $D=0
M340 216 ACTRCLKX 214 VSS N12LL L=6E-08 W=5E-07 $X=21905 $Y=21055 $D=0
M341 216 71 346 VSS N12LL L=6E-08 W=1E-06 $X=21945 $Y=19480 $D=0
M342 106 214 VSS VSS N12LL L=6E-08 W=4E-07 $X=22045 $Y=25095 $D=0
M343 YX[1] 106 58 VSS N12LL L=6E-08 W=1.25E-06 $X=22045 $Y=29015 $D=0
M344 EMCLK 184 218 VSS N12LL L=6E-08 W=1E-06 $X=22060 $Y=12200 $D=0
M345 58 49 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=22155 $Y=3590 $D=0
M346 219 YA[0] 347 VSS N12LL L=6E-08 W=4E-07 $X=22155 $Y=15140 $D=0
M347 214 ACTRCLKX 216 VSS N12LL L=6E-08 W=5E-07 $X=22175 $Y=21055 $D=0
M348 RWLR 215 VSS VSS N12LL L=6E-08 W=1E-06 $X=22310 $Y=33805 $D=0
M349 VSS 215 RWLR VSS N12LL L=6E-08 W=1E-06 $X=22310 $Y=34075 $D=0
M350 218 184 EMCLK VSS N12LL L=6E-08 W=1E-06 $X=22330 $Y=12200 $D=0
M351 VSS 214 106 VSS N12LL L=6E-08 W=4E-07 $X=22335 $Y=25095 $D=0
M352 58 106 YX[1] VSS N12LL L=6E-08 W=1.25E-06 $X=22335 $Y=29015 $D=0
M353 223 217 VSS VSS N12LL L=2E-07 W=4E-07 $X=22385 $Y=1805 $D=0
M354 VSS 49 58 VSS N12LL L=6E-08 W=2.5E-06 $X=22425 $Y=3590 $D=0
M355 108 222 VSS VSS N12LL L=6E-08 W=4E-07 $X=22625 $Y=25095 $D=0
M356 YX[7] 108 58 VSS N12LL L=6E-08 W=1.25E-06 $X=22625 $Y=29015 $D=0
M357 VSS 221 218 VSS N12LL L=6E-08 W=7E-07 $X=22645 $Y=12200 $D=0
M358 58 49 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=22695 $Y=3590 $D=0
M359 71 219 VSS VSS N12LL L=6E-08 W=5E-07 $X=22785 $Y=15060 $D=0
M360 107 ACTRCLKX 222 VSS N12LL L=6E-08 W=5E-07 $X=22785 $Y=21055 $D=0
M361 VSS 108 222 VSS N12LL L=6E-07 W=1.2E-07 $X=22875 $Y=26265 $D=0
M362 221 103 VSS VSS N12LL L=6E-08 W=7E-07 $X=22915 $Y=12200 $D=0
M363 VSS 222 108 VSS N12LL L=6E-08 W=4E-07 $X=22915 $Y=25095 $D=0
M364 58 108 YX[7] VSS N12LL L=6E-08 W=1.25E-06 $X=22915 $Y=29015 $D=0
M365 VSS 49 58 VSS N12LL L=6E-08 W=2.5E-06 $X=22965 $Y=3590 $D=0
M366 348 71 107 VSS N12LL L=6E-08 W=1E-06 $X=23015 $Y=19480 $D=0
M367 222 ACTRCLKX 107 VSS N12LL L=6E-08 W=5E-07 $X=23055 $Y=21055 $D=0
M368 VSS 219 71 VSS N12LL L=6E-08 W=5E-07 $X=23075 $Y=15060 $D=0
M369 109 49 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=23125 $Y=1795 $D=0
M370 108 222 VSS VSS N12LL L=6E-08 W=4E-07 $X=23205 $Y=25095 $D=0
M371 YX[7] 108 58 VSS N12LL L=6E-08 W=1.25E-06 $X=23205 $Y=29015 $D=0
M372 349 68 348 VSS N12LL L=6E-08 W=1E-06 $X=23255 $Y=19480 $D=0
M373 107 ACTRCLKX 222 VSS N12LL L=6E-08 W=5E-07 $X=23335 $Y=21055 $D=0
M374 67 71 VSS VSS N12LL L=6E-08 W=5E-07 $X=23365 $Y=15060 $D=0
M375 VSS 223 109 VSS N12LL L=6E-08 W=7.5E-07 $X=23395 $Y=1795 $D=0
M376 VSS 226 349 VSS N12LL L=6E-08 W=1E-06 $X=23495 $Y=19480 $D=0
M377 VSS 222 108 VSS N12LL L=6E-08 W=4E-07 $X=23495 $Y=25095 $D=0
M378 58 108 YX[7] VSS N12LL L=6E-08 W=1.25E-06 $X=23495 $Y=29015 $D=0
M379 VSS 71 67 VSS N12LL L=6E-08 W=5E-07 $X=23635 $Y=15060 $D=0
M380 109 223 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=23665 $Y=1795 $D=0
M381 350 226 VSS VSS N12LL L=6E-08 W=1E-06 $X=23785 $Y=19480 $D=0
M382 111 224 VSS VSS N12LL L=6E-08 W=4E-07 $X=23785 $Y=25095 $D=0
M383 YX[6] 111 58 VSS N12LL L=6E-08 W=1.25E-06 $X=23785 $Y=29015 $D=0
M384 224 111 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=23865 $Y=26265 $D=0
M385 SACK1 49 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=23925 $Y=10275 $D=0
M386 VSS 49 109 VSS N12LL L=6E-08 W=7.5E-07 $X=23935 $Y=1795 $D=0
M387 224 ACTRCLKX 110 VSS N12LL L=6E-08 W=5E-07 $X=23945 $Y=21055 $D=0
M388 351 68 350 VSS N12LL L=6E-08 W=1E-06 $X=24025 $Y=19480 $D=0
M389 VSS 224 111 VSS N12LL L=6E-08 W=4E-07 $X=24075 $Y=25095 $D=0
M390 58 111 YX[6] VSS N12LL L=6E-08 W=1.25E-06 $X=24075 $Y=29015 $D=0
M391 VSS 49 SACK1 VSS N12LL L=6E-08 W=2.5E-06 $X=24195 $Y=10275 $D=0
M392 110 ACTRCLKX 224 VSS N12LL L=6E-08 W=5E-07 $X=24225 $Y=21055 $D=0
M393 110 67 351 VSS N12LL L=6E-08 W=1E-06 $X=24265 $Y=19480 $D=0
M394 111 224 VSS VSS N12LL L=6E-08 W=4E-07 $X=24365 $Y=25095 $D=0
M395 YX[6] 111 58 VSS N12LL L=6E-08 W=1.25E-06 $X=24365 $Y=29015 $D=0
M396 SACK4 109 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=24465 $Y=10275 $D=0
M397 224 ACTRCLKX 110 VSS N12LL L=6E-08 W=5E-07 $X=24495 $Y=21055 $D=0
M398 228 220 VSS VSS N12LL L=6E-08 W=1.25E-06 $X=24545 $Y=1795 $D=0
M399 VSS 224 111 VSS N12LL L=6E-08 W=4E-07 $X=24655 $Y=25095 $D=0
M400 58 111 YX[6] VSS N12LL L=6E-08 W=1.25E-06 $X=24655 $Y=29015 $D=0
M401 VSS 109 SACK4 VSS N12LL L=6E-08 W=2.5E-06 $X=24735 $Y=10275 $D=0
M402 VSS 49 228 VSS N12LL L=6E-08 W=1.25E-06 $X=24815 $Y=1795 $D=0
M403 352 VDD VSS VSS N12LL L=3E-07 W=4E-07 $X=24865 $Y=15140 $D=0
M404 112 225 VSS VSS N12LL L=6E-08 W=4E-07 $X=24945 $Y=25095 $D=0
M405 YX[4] 112 58 VSS N12LL L=6E-08 W=1.25E-06 $X=24945 $Y=29015 $D=0
M406 DCTRCLK 228 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=25005 $Y=10275 $D=0
M407 228 49 VSS VSS N12LL L=6E-08 W=1.25E-06 $X=25085 $Y=1795 $D=0
M408 113 ACTRCLKX 225 VSS N12LL L=6E-08 W=5E-07 $X=25105 $Y=21055 $D=0
M409 VSS 112 225 VSS N12LL L=6E-07 W=1.2E-07 $X=25195 $Y=26265 $D=0
M410 VSS 225 112 VSS N12LL L=6E-08 W=4E-07 $X=25235 $Y=25095 $D=0
M411 58 112 YX[4] VSS N12LL L=6E-08 W=1.25E-06 $X=25235 $Y=29015 $D=0
M412 VSS 228 DCTRCLK VSS N12LL L=6E-08 W=2.5E-06 $X=25275 $Y=10275 $D=0
M413 227 YA[1] 352 VSS N12LL L=6E-08 W=4E-07 $X=25335 $Y=15140 $D=0
M414 353 67 113 VSS N12LL L=6E-08 W=1E-06 $X=25335 $Y=19480 $D=0
M415 VSS 220 228 VSS N12LL L=6E-08 W=1.25E-06 $X=25355 $Y=1795 $D=0
M416 225 ACTRCLKX 113 VSS N12LL L=6E-08 W=5E-07 $X=25375 $Y=21055 $D=0
M417 112 225 VSS VSS N12LL L=6E-08 W=4E-07 $X=25525 $Y=25095 $D=0
M418 YX[4] 112 58 VSS N12LL L=6E-08 W=1.25E-06 $X=25525 $Y=29015 $D=0
M419 ACTRCLK 228 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=25545 $Y=10275 $D=0
M420 354 230 353 VSS N12LL L=6E-08 W=1E-06 $X=25575 $Y=19480 $D=0
M421 113 ACTRCLKX 225 VSS N12LL L=6E-08 W=5E-07 $X=25655 $Y=21055 $D=0
M422 VSS 228 ACTRCLK VSS N12LL L=6E-08 W=2.5E-06 $X=25815 $Y=10275 $D=0
M423 VSS 226 354 VSS N12LL L=6E-08 W=1E-06 $X=25815 $Y=19480 $D=0
M424 VSS 225 112 VSS N12LL L=6E-08 W=4E-07 $X=25815 $Y=25095 $D=0
M425 58 112 YX[4] VSS N12LL L=6E-08 W=1.25E-06 $X=25815 $Y=29015 $D=0
M426 231 228 VSS VSS N12LL L=6E-08 W=1E-06 $X=25945 $Y=1795 $D=0
M427 68 227 VSS VSS N12LL L=6E-08 W=5E-07 $X=25965 $Y=15060 $D=0
M428 ACTRCLKX ACTRCLK VSS VSS N12LL L=6E-08 W=2.5E-06 $X=26085 $Y=10275 $D=0
M429 355 226 VSS VSS N12LL L=6E-08 W=1E-06 $X=26105 $Y=19480 $D=0
M430 114 229 VSS VSS N12LL L=6E-08 W=4E-07 $X=26105 $Y=25095 $D=0
M431 YX[5] 114 58 VSS N12LL L=6E-08 W=1.25E-06 $X=26105 $Y=29015 $D=0
M432 229 114 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=26185 $Y=26265 $D=0
M433 VSS 228 231 VSS N12LL L=6E-08 W=1E-06 $X=26215 $Y=1795 $D=0
M434 VSS 227 68 VSS N12LL L=6E-08 W=5E-07 $X=26255 $Y=15060 $D=0
M435 229 ACTRCLKX 232 VSS N12LL L=6E-08 W=5E-07 $X=26265 $Y=21055 $D=0
M436 356 230 355 VSS N12LL L=6E-08 W=1E-06 $X=26345 $Y=19480 $D=0
M437 VSS ACTRCLK ACTRCLKX VSS N12LL L=6E-08 W=2.5E-06 $X=26355 $Y=10275 $D=0
M438 VSS 229 114 VSS N12LL L=6E-08 W=4E-07 $X=26395 $Y=25095 $D=0
M439 58 114 YX[5] VSS N12LL L=6E-08 W=1.25E-06 $X=26395 $Y=29015 $D=0
M440 231 228 VSS VSS N12LL L=6E-08 W=1E-06 $X=26485 $Y=1795 $D=0
M441 230 68 VSS VSS N12LL L=6E-08 W=5E-07 $X=26545 $Y=15060 $D=0
M442 232 ACTRCLKX 229 VSS N12LL L=6E-08 W=5E-07 $X=26545 $Y=21055 $D=0
M443 232 71 356 VSS N12LL L=6E-08 W=1E-06 $X=26585 $Y=19480 $D=0
M444 DCTRCLKX 231 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=26625 $Y=10275 $D=0
M445 114 229 VSS VSS N12LL L=6E-08 W=4E-07 $X=26685 $Y=25095 $D=0
M446 YX[5] 114 58 VSS N12LL L=6E-08 W=1.25E-06 $X=26685 $Y=29015 $D=0
M447 VSS 68 230 VSS N12LL L=6E-08 W=5E-07 $X=26815 $Y=15060 $D=0
M448 229 ACTRCLKX 232 VSS N12LL L=6E-08 W=5E-07 $X=26815 $Y=21055 $D=0
M449 VSS 231 DCTRCLKX VSS N12LL L=6E-08 W=2.5E-06 $X=26895 $Y=10275 $D=0
M450 VSS 229 114 VSS N12LL L=6E-08 W=4E-07 $X=26975 $Y=25095 $D=0
M451 58 114 YX[5] VSS N12LL L=6E-08 W=1.25E-06 $X=26975 $Y=29015 $D=0
M452 357 XA[3] 123 VDD P12LL L=6E-08 W=4E-07 $X=640 $Y=2130 $D=2
M453 VDD RDE 357 VDD P12LL L=6E-08 W=4E-07 $X=910 $Y=2130 $D=2
M454 RWLL 131 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=940 $Y=33805 $D=2
M455 VDD 131 RWLL VDD P12LL L=6E-08 W=2.5E-06 $X=940 $Y=34075 $D=2
M456 124 123 VDD VDD P12LL L=3E-07 W=4E-07 $X=1220 $Y=2130 $D=2
M457 VDD 124 125 VDD P12LL L=6E-08 W=4E-07 $X=2080 $Y=2130 $D=2
M458 127 125 VDD VDD P12LL L=6E-08 W=2E-06 $X=2400 $Y=530 $D=2
M459 VDD ZAX 128 VDD P12LL L=3E-07 W=1.2E-07 $X=3070 $Y=195 $D=2
M460 127 ACTRCLK 128 VDD P12LL L=6E-08 W=1.245E-06 $X=3115 $Y=1285 $D=2
M461 128 ACTRCLK 127 VDD P12LL L=6E-08 W=1.245E-06 $X=3385 $Y=1285 $D=2
M462 ZAX 128 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=3995 $Y=5 $D=2
M463 VDD 128 ZAX VDD P12LL L=6E-08 W=2.5E-06 $X=4265 $Y=5 $D=2
M464 ZAX 128 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=4535 $Y=5 $D=2
M465 VDD 128 ZAX VDD P12LL L=6E-08 W=2.5E-06 $X=4805 $Y=5 $D=2
M466 PXA[3] 132 VDD VDD P12LL L=6E-08 W=3.5E-06 $X=5015 $Y=27075 $D=2
M467 130 142 VDD VDD P12LL L=6E-08 W=1.5E-06 $X=5035 $Y=15400 $D=2
M468 358 134 142 VDD P12LL L=6E-08 W=7E-07 $X=5095 $Y=10320 $D=2
M469 133 128 VDD VDD P12LL L=6E-08 W=2E-06 $X=5115 $Y=505 $D=2
M470 132 ACTRCLK 130 VDD P12LL L=6E-08 W=2.5E-06 $X=5160 $Y=20435 $D=2
M471 136 PXA[2] VDD VDD P12LL L=3E-07 W=1.2E-07 $X=5295 $Y=31225 $D=2
M472 VDD 132 PXA[3] VDD P12LL L=6E-08 W=3.5E-06 $X=5305 $Y=27075 $D=2
M473 VDD 140 130 VDD P12LL L=6E-08 W=1.5E-06 $X=5320 $Y=15400 $D=2
M474 VDD RDE 358 VDD P12LL L=6E-08 W=7E-07 $X=5385 $Y=10320 $D=2
M475 VDD XA[3] 134 VDD P12LL L=6E-08 W=4E-07 $X=5440 $Y=8705 $D=2
M476 VDD PXA[3] 132 VDD P12LL L=3E-07 W=1.2E-07 $X=5550 $Y=31880 $D=2
M477 135 140 VDD VDD P12LL L=6E-08 W=1.5E-06 $X=5580 $Y=15400 $D=2
M478 PXA[2] 136 VDD VDD P12LL L=6E-08 W=3.5E-06 $X=5595 $Y=27075 $D=2
M479 359 RDE VDD VDD P12LL L=6E-08 W=1.4E-06 $X=5675 $Y=9620 $D=2
M480 ZA 133 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=5735 $Y=5 $D=2
M481 135 ACTRCLK 136 VDD P12LL L=6E-08 W=2.5E-06 $X=5740 $Y=20435 $D=2
M482 137 134 VDD VDD P12LL L=6E-08 W=4E-07 $X=5765 $Y=8705 $D=2
M483 VDD 73 135 VDD P12LL L=6E-08 W=1.5E-06 $X=5865 $Y=15400 $D=2
M484 VDD 136 PXA[2] VDD P12LL L=6E-08 W=3.5E-06 $X=5885 $Y=27075 $D=2
M485 73 137 359 VDD P12LL L=6E-08 W=1.4E-06 $X=5965 $Y=9620 $D=2
M486 VDD 133 ZA VDD P12LL L=6E-08 W=2.5E-06 $X=6005 $Y=5 $D=2
M487 PXA[0] 138 VDD VDD P12LL L=6E-08 W=3.5E-06 $X=6225 $Y=27075 $D=2
M488 139 73 VDD VDD P12LL L=6E-08 W=1.5E-06 $X=6245 $Y=15400 $D=2
M489 ZA 133 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=6275 $Y=5 $D=2
M490 141 PXA[1] VDD VDD P12LL L=3E-07 W=1.2E-07 $X=6320 $Y=31880 $D=2
M491 138 ACTRCLK 139 VDD P12LL L=6E-08 W=2.5E-06 $X=6370 $Y=20435 $D=2
M492 VDD 138 PXA[0] VDD P12LL L=6E-08 W=3.5E-06 $X=6515 $Y=27075 $D=2
M493 VDD 145 139 VDD P12LL L=6E-08 W=1.5E-06 $X=6530 $Y=15400 $D=2
M494 VDD 133 ZA VDD P12LL L=6E-08 W=2.5E-06 $X=6545 $Y=5 $D=2
M495 VDD PXA[0] 138 VDD P12LL L=3E-07 W=1.2E-07 $X=6575 $Y=31225 $D=2
M496 360 VSS VDD VDD P12LL L=1E-07 W=4E-07 $X=6700 $Y=8705 $D=2
M497 143 145 VDD VDD P12LL L=6E-08 W=1.5E-06 $X=6790 $Y=15400 $D=2
M498 PXA[1] 141 VDD VDD P12LL L=6E-08 W=3.5E-06 $X=6805 $Y=27075 $D=2
M499 VDD 144 140 VDD P12LL L=6E-08 W=1.4E-06 $X=6820 $Y=9620 $D=2
M500 143 ACTRCLK 141 VDD P12LL L=6E-08 W=2.5E-06 $X=6950 $Y=20435 $D=2
M501 144 XA[4] 360 VDD P12LL L=6E-08 W=4E-07 $X=7000 $Y=8705 $D=2
M502 131 209 VDD VDD P12LL L=6E-08 W=1E-06 $X=7070 $Y=33805 $D=2
M503 VDD 209 131 VDD P12LL L=6E-08 W=1E-06 $X=7070 $Y=34075 $D=2
M504 VDD 142 143 VDD P12LL L=6E-08 W=1.5E-06 $X=7075 $Y=15400 $D=2
M505 VDD 141 PXA[1] VDD P12LL L=6E-08 W=3.5E-06 $X=7095 $Y=27075 $D=2
M506 145 140 VDD VDD P12LL L=6E-08 W=1.4E-06 $X=7110 $Y=9620 $D=2
M507 131 198 58 VDD P12LL L=6E-08 W=5E-07 $X=8570 $Y=33805 $D=2
M508 58 198 131 VDD P12LL L=6E-08 W=5E-07 $X=8570 $Y=34075 $D=2
M509 76 149 VDD VDD P12LL L=6E-08 W=4E-07 $X=8705 $Y=24010 $D=2
M510 FCKX[3] 149 58 VDD P12LL L=6E-08 W=1.25E-06 $X=8705 $Y=27205 $D=2
M511 FCKX[3] 76 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=8705 $Y=30765 $D=2
M512 161 188 VDD VDD P12LL L=6E-08 W=1E-06 $X=8865 $Y=16080 $D=2
M513 152 ACTRCLK 149 VDD P12LL L=6E-08 W=5E-07 $X=8865 $Y=22055 $D=2
M514 VDD 61 152 VDD P12LL L=6E-08 W=1E-06 $X=8995 $Y=17910 $D=2
M515 VDD 149 76 VDD P12LL L=6E-08 W=4E-07 $X=8995 $Y=24010 $D=2
M516 58 149 FCKX[3] VDD P12LL L=6E-08 W=1.25E-06 $X=8995 $Y=27205 $D=2
M517 VDD 76 FCKX[3] VDD P12LL L=6E-08 W=1.25E-06 $X=8995 $Y=30765 $D=2
M518 VDD 188 161 VDD P12LL L=6E-08 W=1E-06 $X=9135 $Y=16080 $D=2
M519 149 ACTRCLK 152 VDD P12LL L=6E-08 W=5E-07 $X=9135 $Y=22055 $D=2
M520 VDD 76 149 VDD P12LL L=3E-07 W=1.2E-07 $X=9245 $Y=23170 $D=2
M521 152 60 VDD VDD P12LL L=6E-08 W=1E-06 $X=9285 $Y=17910 $D=2
M522 76 149 VDD VDD P12LL L=6E-08 W=4E-07 $X=9285 $Y=24010 $D=2
M523 FCKX[3] 149 58 VDD P12LL L=6E-08 W=1.25E-06 $X=9285 $Y=27205 $D=2
M524 FCKX[3] 76 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=9285 $Y=30765 $D=2
M525 152 ACTRCLK 149 VDD P12LL L=6E-08 W=5E-07 $X=9415 $Y=22055 $D=2
M526 188 155 VDD VDD P12LL L=6E-08 W=1E-06 $X=9425 $Y=16080 $D=2
M527 VDD 161 152 VDD P12LL L=6E-08 W=1E-06 $X=9575 $Y=17910 $D=2
M528 VDD 149 76 VDD P12LL L=6E-08 W=4E-07 $X=9575 $Y=24010 $D=2
M529 58 149 FCKX[3] VDD P12LL L=6E-08 W=1.25E-06 $X=9575 $Y=27205 $D=2
M530 VDD 76 FCKX[3] VDD P12LL L=6E-08 W=1.25E-06 $X=9575 $Y=30765 $D=2
M531 VDD 155 188 VDD P12LL L=6E-08 W=1E-06 $X=9715 $Y=16080 $D=2
M532 78 161 VDD VDD P12LL L=6E-08 W=1E-06 $X=9865 $Y=17910 $D=2
M533 80 156 VDD VDD P12LL L=6E-08 W=4E-07 $X=9865 $Y=24010 $D=2
M534 FCKX[2] 156 58 VDD P12LL L=6E-08 W=1.25E-06 $X=9865 $Y=27205 $D=2
M535 FCKX[2] 80 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=9865 $Y=30765 $D=2
M536 156 80 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=9955 $Y=23170 $D=2
M537 156 ACTRCLK 78 VDD P12LL L=6E-08 W=5E-07 $X=10025 $Y=22055 $D=2
M538 VDD 60 78 VDD P12LL L=6E-08 W=1E-06 $X=10155 $Y=17910 $D=2
M539 VDD 156 80 VDD P12LL L=6E-08 W=4E-07 $X=10155 $Y=24010 $D=2
M540 58 156 FCKX[2] VDD P12LL L=6E-08 W=1.25E-06 $X=10155 $Y=27205 $D=2
M541 VDD 80 FCKX[2] VDD P12LL L=6E-08 W=1.25E-06 $X=10155 $Y=30765 $D=2
M542 78 ACTRCLK 156 VDD P12LL L=6E-08 W=5E-07 $X=10305 $Y=22055 $D=2
M543 361 XA[2] 155 VDD P12LL L=6E-08 W=4E-07 $X=10345 $Y=16410 $D=2
M544 78 59 VDD VDD P12LL L=6E-08 W=1E-06 $X=10445 $Y=17910 $D=2
M545 80 156 VDD VDD P12LL L=6E-08 W=4E-07 $X=10445 $Y=24010 $D=2
M546 FCKX[2] 156 58 VDD P12LL L=6E-08 W=1.25E-06 $X=10445 $Y=27205 $D=2
M547 FCKX[2] 80 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=10445 $Y=30765 $D=2
M548 156 ACTRCLK 78 VDD P12LL L=6E-08 W=5E-07 $X=10575 $Y=22055 $D=2
M549 VDD VSS 361 VDD P12LL L=1E-07 W=4E-07 $X=10635 $Y=16410 $D=2
M550 VDD 156 80 VDD P12LL L=6E-08 W=4E-07 $X=10735 $Y=24010 $D=2
M551 58 156 FCKX[2] VDD P12LL L=6E-08 W=1.25E-06 $X=10735 $Y=27205 $D=2
M552 VDD 80 FCKX[2] VDD P12LL L=6E-08 W=1.25E-06 $X=10735 $Y=30765 $D=2
M553 82 160 VDD VDD P12LL L=6E-08 W=4E-07 $X=11025 $Y=24010 $D=2
M554 FCKX[0] 160 58 VDD P12LL L=6E-08 W=1.25E-06 $X=11025 $Y=27205 $D=2
M555 FCKX[0] 82 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=11025 $Y=30765 $D=2
M556 84 ACTRCLK 160 VDD P12LL L=6E-08 W=5E-07 $X=11185 $Y=22055 $D=2
M557 VDD 59 84 VDD P12LL L=6E-08 W=1E-06 $X=11315 $Y=17910 $D=2
M558 VDD 160 82 VDD P12LL L=6E-08 W=4E-07 $X=11315 $Y=24010 $D=2
M559 58 160 FCKX[0] VDD P12LL L=6E-08 W=1.25E-06 $X=11315 $Y=27205 $D=2
M560 VDD 82 FCKX[0] VDD P12LL L=6E-08 W=1.25E-06 $X=11315 $Y=30765 $D=2
M561 160 ACTRCLK 84 VDD P12LL L=6E-08 W=5E-07 $X=11455 $Y=22055 $D=2
M562 VDD 82 160 VDD P12LL L=3E-07 W=1.2E-07 $X=11565 $Y=23170 $D=2
M563 84 194 VDD VDD P12LL L=6E-08 W=1E-06 $X=11605 $Y=17910 $D=2
M564 82 160 VDD VDD P12LL L=6E-08 W=4E-07 $X=11605 $Y=24010 $D=2
M565 FCKX[0] 160 58 VDD P12LL L=6E-08 W=1.25E-06 $X=11605 $Y=27205 $D=2
M566 FCKX[0] 82 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=11605 $Y=30765 $D=2
M567 83 162 VDD VDD P12LL L=6E-08 W=4E-07 $X=11690 $Y=13290 $D=2
M568 84 ACTRCLK 160 VDD P12LL L=6E-08 W=5E-07 $X=11735 $Y=22055 $D=2
M569 VDD S[0] 162 VDD P12LL L=6E-08 W=4E-07 $X=11790 $Y=9890 $D=2
M570 VDD 161 84 VDD P12LL L=6E-08 W=1E-06 $X=11895 $Y=17910 $D=2
M571 VDD 160 82 VDD P12LL L=6E-08 W=4E-07 $X=11895 $Y=24010 $D=2
M572 58 160 FCKX[0] VDD P12LL L=6E-08 W=1.25E-06 $X=11895 $Y=27205 $D=2
M573 VDD 82 FCKX[0] VDD P12LL L=6E-08 W=1.25E-06 $X=11895 $Y=30765 $D=2
M574 VDD 85 163 VDD P12LL L=3E-07 W=1.2E-07 $X=11945 $Y=8760 $D=2
M575 VDD 88 83 VDD P12LL L=6E-08 W=4E-07 $X=11960 $Y=13290 $D=2
M576 164 WEN VDD VDD P12LL L=6E-08 W=4E-07 $X=11990 $Y=475 $D=2
M577 173 162 VDD VDD P12LL L=6E-08 W=4E-07 $X=12060 $Y=9890 $D=2
M578 166 161 VDD VDD P12LL L=6E-08 W=1E-06 $X=12185 $Y=17910 $D=2
M579 86 165 VDD VDD P12LL L=6E-08 W=4E-07 $X=12185 $Y=24010 $D=2
M580 FCKX[1] 165 58 VDD P12LL L=6E-08 W=1.25E-06 $X=12185 $Y=27205 $D=2
M581 FCKX[1] 86 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=12185 $Y=30765 $D=2
M582 208 83 VDD VDD P12LL L=6E-08 W=4E-07 $X=12230 $Y=13290 $D=2
M583 165 86 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=12275 $Y=23170 $D=2
M584 VDD 163 85 VDD P12LL L=6E-08 W=1E-06 $X=12325 $Y=6710 $D=2
M585 165 ACTRCLK 166 VDD P12LL L=6E-08 W=5E-07 $X=12345 $Y=22055 $D=2
M586 VDD 194 166 VDD P12LL L=6E-08 W=1E-06 $X=12475 $Y=17910 $D=2
M587 VDD 165 86 VDD P12LL L=6E-08 W=4E-07 $X=12475 $Y=24010 $D=2
M588 58 165 FCKX[1] VDD P12LL L=6E-08 W=1.25E-06 $X=12475 $Y=27205 $D=2
M589 VDD 86 FCKX[1] VDD P12LL L=6E-08 W=1.25E-06 $X=12475 $Y=30765 $D=2
M590 363 VSS VDD VDD P12LL L=1E-07 W=4E-07 $X=12545 $Y=16410 $D=2
M591 168 85 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=12625 $Y=6710 $D=2
M592 166 ACTRCLK 165 VDD P12LL L=6E-08 W=5E-07 $X=12625 $Y=22055 $D=2
M593 VDD 164 167 VDD P12LL L=3E-07 W=4E-07 $X=12695 $Y=475 $D=2
M594 166 61 VDD VDD P12LL L=6E-08 W=1E-06 $X=12765 $Y=17910 $D=2
M595 86 165 VDD VDD P12LL L=6E-08 W=4E-07 $X=12765 $Y=24010 $D=2
M596 FCKX[1] 165 58 VDD P12LL L=6E-08 W=1.25E-06 $X=12765 $Y=27205 $D=2
M597 FCKX[1] 86 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=12765 $Y=30765 $D=2
M598 VDD 49 168 VDD P12LL L=6E-08 W=2.5E-06 $X=12875 $Y=6710 $D=2
M599 169 XA[0] 363 VDD P12LL L=6E-08 W=4E-07 $X=12875 $Y=16410 $D=2
M600 165 ACTRCLK 166 VDD P12LL L=6E-08 W=5E-07 $X=12895 $Y=22055 $D=2
M601 87 173 VDD VDD P12LL L=6E-08 W=4E-07 $X=12920 $Y=13290 $D=2
M602 VDD 165 86 VDD P12LL L=6E-08 W=4E-07 $X=13055 $Y=24010 $D=2
M603 58 165 FCKX[1] VDD P12LL L=6E-08 W=1.25E-06 $X=13055 $Y=27205 $D=2
M604 VDD 86 FCKX[1] VDD P12LL L=6E-08 W=1.25E-06 $X=13055 $Y=30765 $D=2
M605 WE 168 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=13125 $Y=6710 $D=2
M606 VDD 174 87 VDD P12LL L=6E-08 W=4E-07 $X=13260 $Y=13290 $D=2
M607 171 167 VDD VDD P12LL L=2E-07 W=4E-07 $X=13325 $Y=475 $D=2
M608 89 170 VDD VDD P12LL L=6E-08 W=4E-07 $X=13345 $Y=24010 $D=2
M609 FCKX[7] 170 58 VDD P12LL L=6E-08 W=1.25E-06 $X=13345 $Y=27205 $D=2
M610 FCKX[7] 89 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=13345 $Y=30765 $D=2
M611 VDD 168 WE VDD P12LL L=6E-08 W=2.5E-06 $X=13375 $Y=6710 $D=2
M612 VDD S[1] 174 VDD P12LL L=6E-08 W=4E-07 $X=13405 $Y=9890 $D=2
M613 61 169 VDD VDD P12LL L=6E-08 W=1E-06 $X=13505 $Y=16080 $D=2
M614 90 ACTRCLK 170 VDD P12LL L=6E-08 W=5E-07 $X=13505 $Y=22055 $D=2
M615 172 87 VDD VDD P12LL L=6E-08 W=4E-07 $X=13530 $Y=13290 $D=2
M616 WE 168 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=13625 $Y=6710 $D=2
M617 VDD 61 90 VDD P12LL L=6E-08 W=1E-06 $X=13635 $Y=17910 $D=2
M618 VDD 170 89 VDD P12LL L=6E-08 W=4E-07 $X=13635 $Y=24010 $D=2
M619 58 170 FCKX[7] VDD P12LL L=6E-08 W=1.25E-06 $X=13635 $Y=27205 $D=2
M620 VDD 89 FCKX[7] VDD P12LL L=6E-08 W=1.25E-06 $X=13635 $Y=30765 $D=2
M621 88 174 VDD VDD P12LL L=6E-08 W=4E-07 $X=13665 $Y=9890 $D=2
M622 170 ACTRCLK 90 VDD P12LL L=6E-08 W=5E-07 $X=13775 $Y=22055 $D=2
M623 VDD 169 61 VDD P12LL L=6E-08 W=1E-06 $X=13795 $Y=16080 $D=2
M624 VDD 168 WE VDD P12LL L=6E-08 W=2.5E-06 $X=13875 $Y=6710 $D=2
M625 VDD 89 170 VDD P12LL L=3E-07 W=1.2E-07 $X=13885 $Y=23170 $D=2
M626 90 60 VDD VDD P12LL L=6E-08 W=1E-06 $X=13925 $Y=17910 $D=2
M627 89 170 VDD VDD P12LL L=6E-08 W=4E-07 $X=13925 $Y=24010 $D=2
M628 FCKX[7] 170 58 VDD P12LL L=6E-08 W=1.25E-06 $X=13925 $Y=27205 $D=2
M629 FCKX[7] 89 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=13925 $Y=30765 $D=2
M630 90 ACTRCLK 170 VDD P12LL L=6E-08 W=5E-07 $X=14055 $Y=22055 $D=2
M631 59 61 VDD VDD P12LL L=6E-08 W=1E-06 $X=14085 $Y=16080 $D=2
M632 175 171 VDD VDD P12LL L=6E-08 W=1E-06 $X=14105 $Y=-50 $D=2
M633 181 162 VDD VDD P12LL L=6E-08 W=4E-07 $X=14130 $Y=13290 $D=2
M634 VDD 188 90 VDD P12LL L=6E-08 W=1E-06 $X=14215 $Y=17910 $D=2
M635 VDD 170 89 VDD P12LL L=6E-08 W=4E-07 $X=14215 $Y=24010 $D=2
M636 58 170 FCKX[7] VDD P12LL L=6E-08 W=1.25E-06 $X=14215 $Y=27205 $D=2
M637 VDD 89 FCKX[7] VDD P12LL L=6E-08 W=1.25E-06 $X=14215 $Y=30765 $D=2
M638 VDD 185 198 VDD P12LL L=6E-08 W=8E-07 $X=14240 $Y=34560 $D=2
M639 209 198 VDD VDD P12LL L=6E-08 W=8E-07 $X=14240 $Y=34830 $D=2
M640 183 173 VDD VDD P12LL L=6E-08 W=4E-07 $X=14260 $Y=9890 $D=2
M641 VDD RDE 182 VDD P12LL L=6E-08 W=8E-07 $X=14300 $Y=33350 $D=2
M642 176 182 VDD VDD P12LL L=6E-08 W=8E-07 $X=14300 $Y=33620 $D=2
M643 185 ACTRCLK 176 VDD P12LL L=6E-08 W=1E-06 $X=14300 $Y=33930 $D=2
M644 VDD 61 59 VDD P12LL L=6E-08 W=1E-06 $X=14355 $Y=16080 $D=2
M645 163 ACTRCLK 175 VDD P12LL L=6E-08 W=1E-06 $X=14375 $Y=-50 $D=2
M646 VDD 174 181 VDD P12LL L=6E-08 W=4E-07 $X=14400 $Y=13290 $D=2
M647 VDD 177 196 VDD P12LL L=6E-08 W=2.5E-06 $X=14415 $Y=6790 $D=2
M648 91 188 VDD VDD P12LL L=6E-08 W=1E-06 $X=14505 $Y=17910 $D=2
M649 92 180 VDD VDD P12LL L=6E-08 W=4E-07 $X=14505 $Y=24010 $D=2
M650 FCKX[6] 180 58 VDD P12LL L=6E-08 W=1.25E-06 $X=14505 $Y=27205 $D=2
M651 FCKX[6] 92 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=14505 $Y=30765 $D=2
M652 VDD 88 183 VDD P12LL L=6E-08 W=4E-07 $X=14530 $Y=9890 $D=2
M653 180 92 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=14595 $Y=23170 $D=2
M654 180 ACTRCLK 91 VDD P12LL L=6E-08 W=5E-07 $X=14665 $Y=22055 $D=2
M655 178 181 VDD VDD P12LL L=6E-08 W=4E-07 $X=14670 $Y=13290 $D=2
M656 177 FB VDD VDD P12LL L=6E-08 W=8E-07 $X=14745 $Y=6790 $D=2
M657 VDD 60 91 VDD P12LL L=6E-08 W=1E-06 $X=14795 $Y=17910 $D=2
M658 VDD 180 92 VDD P12LL L=6E-08 W=4E-07 $X=14795 $Y=24010 $D=2
M659 58 180 FCKX[6] VDD P12LL L=6E-08 W=1.25E-06 $X=14795 $Y=27205 $D=2
M660 VDD 92 FCKX[6] VDD P12LL L=6E-08 W=1.25E-06 $X=14795 $Y=30765 $D=2
M661 184 183 VDD VDD P12LL L=6E-08 W=4E-07 $X=14800 $Y=9890 $D=2
M662 91 ACTRCLK 180 VDD P12LL L=6E-08 W=5E-07 $X=14945 $Y=22055 $D=2
M663 VDD CLK 179 VDD P12LL L=6E-08 W=4E-07 $X=14955 $Y=500 $D=2
M664 91 59 VDD VDD P12LL L=6E-08 W=1E-06 $X=15085 $Y=17910 $D=2
M665 92 180 VDD VDD P12LL L=6E-08 W=4E-07 $X=15085 $Y=24010 $D=2
M666 FCKX[6] 180 58 VDD P12LL L=6E-08 W=1.25E-06 $X=15085 $Y=27205 $D=2
M667 FCKX[6] 92 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=15085 $Y=30765 $D=2
M668 180 ACTRCLK 91 VDD P12LL L=6E-08 W=5E-07 $X=15215 $Y=22055 $D=2
M669 364 CLK VDD VDD P12LL L=6E-08 W=1E-06 $X=15310 $Y=-100 $D=2
M670 VDD 180 92 VDD P12LL L=6E-08 W=4E-07 $X=15375 $Y=24010 $D=2
M671 58 180 FCKX[6] VDD P12LL L=6E-08 W=1.25E-06 $X=15375 $Y=27205 $D=2
M672 VDD 92 FCKX[6] VDD P12LL L=6E-08 W=1.25E-06 $X=15375 $Y=30765 $D=2
M673 190 CEN 364 VDD P12LL L=6E-08 W=1E-06 $X=15545 $Y=-100 $D=2
M674 93 186 VDD VDD P12LL L=6E-08 W=4E-07 $X=15665 $Y=24010 $D=2
M675 FCKX[4] 186 58 VDD P12LL L=6E-08 W=1.25E-06 $X=15665 $Y=27205 $D=2
M676 FCKX[4] 93 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=15665 $Y=30765 $D=2
M677 365 VSS VDD VDD P12LL L=1E-07 W=4E-07 $X=15725 $Y=16410 $D=2
M678 94 ACTRCLK 186 VDD P12LL L=6E-08 W=5E-07 $X=15825 $Y=22055 $D=2
M679 EMCLK 181 187 VDD P12LL L=6E-08 W=1.25E-06 $X=15860 $Y=10100 $D=2
M680 VDD 192 190 VDD P12LL L=3E-07 W=1.2E-07 $X=15905 $Y=780 $D=2
M681 VDD 59 94 VDD P12LL L=6E-08 W=1E-06 $X=15955 $Y=17910 $D=2
M682 VDD 186 93 VDD P12LL L=6E-08 W=4E-07 $X=15955 $Y=24010 $D=2
M683 58 186 FCKX[4] VDD P12LL L=6E-08 W=1.25E-06 $X=15955 $Y=27205 $D=2
M684 VDD 93 FCKX[4] VDD P12LL L=6E-08 W=1.25E-06 $X=15955 $Y=30765 $D=2
M685 189 XA[1] 365 VDD P12LL L=6E-08 W=4E-07 $X=16055 $Y=16410 $D=2
M686 186 ACTRCLK 94 VDD P12LL L=6E-08 W=5E-07 $X=16095 $Y=22055 $D=2
M687 187 181 EMCLK VDD P12LL L=6E-08 W=1.25E-06 $X=16130 $Y=10100 $D=2
M688 VDD 198 185 VDD P12LL L=3E-07 W=1.2E-07 $X=16135 $Y=33865 $D=2
M689 VDD 93 186 VDD P12LL L=3E-07 W=1.2E-07 $X=16205 $Y=23170 $D=2
M690 94 194 VDD VDD P12LL L=6E-08 W=1E-06 $X=16245 $Y=17910 $D=2
M691 93 186 VDD VDD P12LL L=6E-08 W=4E-07 $X=16245 $Y=24010 $D=2
M692 FCKX[4] 186 58 VDD P12LL L=6E-08 W=1.25E-06 $X=16245 $Y=27205 $D=2
M693 FCKX[4] 93 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=16245 $Y=30765 $D=2
M694 94 ACTRCLK 186 VDD P12LL L=6E-08 W=5E-07 $X=16375 $Y=22055 $D=2
M695 VDD 191 187 VDD P12LL L=6E-08 W=1.4E-06 $X=16460 $Y=9950 $D=2
M696 VDD 188 94 VDD P12LL L=6E-08 W=1E-06 $X=16535 $Y=17910 $D=2
M697 VDD 186 93 VDD P12LL L=6E-08 W=4E-07 $X=16535 $Y=24010 $D=2
M698 58 186 FCKX[4] VDD P12LL L=6E-08 W=1.25E-06 $X=16535 $Y=27205 $D=2
M699 VDD 93 FCKX[4] VDD P12LL L=6E-08 W=1.25E-06 $X=16535 $Y=30765 $D=2
M700 60 189 VDD VDD P12LL L=6E-08 W=1E-06 $X=16685 $Y=16080 $D=2
M701 195 188 VDD VDD P12LL L=6E-08 W=1E-06 $X=16825 $Y=17910 $D=2
M702 96 193 VDD VDD P12LL L=6E-08 W=4E-07 $X=16825 $Y=24010 $D=2
M703 FCKX[5] 193 58 VDD P12LL L=6E-08 W=1.25E-06 $X=16825 $Y=27205 $D=2
M704 FCKX[5] 96 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=16825 $Y=30765 $D=2
M705 192 190 VDD VDD P12LL L=6E-08 W=8E-07 $X=16835 $Y=150 $D=2
M706 193 96 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=16915 $Y=23170 $D=2
M707 VDD 189 60 VDD P12LL L=6E-08 W=1E-06 $X=16975 $Y=16080 $D=2
M708 193 ACTRCLK 195 VDD P12LL L=6E-08 W=5E-07 $X=16985 $Y=22055 $D=2
M709 VDD 194 195 VDD P12LL L=6E-08 W=1E-06 $X=17115 $Y=17910 $D=2
M710 VDD 193 96 VDD P12LL L=6E-08 W=4E-07 $X=17115 $Y=24010 $D=2
M711 58 193 FCKX[5] VDD P12LL L=6E-08 W=1.25E-06 $X=17115 $Y=27205 $D=2
M712 VDD 96 FCKX[5] VDD P12LL L=6E-08 W=1.25E-06 $X=17115 $Y=30765 $D=2
M713 VDD 221 FB VDD P12LL L=6E-08 W=2.4E-06 $X=17195 $Y=6890 $D=2
M714 194 60 VDD VDD P12LL L=6E-08 W=1E-06 $X=17265 $Y=16080 $D=2
M715 195 ACTRCLK 193 VDD P12LL L=6E-08 W=5E-07 $X=17265 $Y=22055 $D=2
M716 VDD 203 191 VDD P12LL L=1.5E-07 W=7E-07 $X=17345 $Y=10600 $D=2
M717 195 61 VDD VDD P12LL L=6E-08 W=1E-06 $X=17405 $Y=17910 $D=2
M718 96 193 VDD VDD P12LL L=6E-08 W=4E-07 $X=17405 $Y=24010 $D=2
M719 FCKX[5] 193 58 VDD P12LL L=6E-08 W=1.25E-06 $X=17405 $Y=27205 $D=2
M720 FCKX[5] 96 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=17405 $Y=30765 $D=2
M721 103 196 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=17475 $Y=6890 $D=2
M722 367 192 197 VDD P12LL L=6E-08 W=1E-06 $X=17515 $Y=-100 $D=2
M723 VDD 60 194 VDD P12LL L=6E-08 W=1E-06 $X=17535 $Y=16080 $D=2
M724 193 ACTRCLK 195 VDD P12LL L=6E-08 W=5E-07 $X=17535 $Y=22055 $D=2
M725 VDD 193 96 VDD P12LL L=6E-08 W=4E-07 $X=17695 $Y=24010 $D=2
M726 58 193 FCKX[5] VDD P12LL L=6E-08 W=1.25E-06 $X=17695 $Y=27205 $D=2
M727 VDD 96 FCKX[5] VDD P12LL L=6E-08 W=1.25E-06 $X=17695 $Y=30765 $D=2
M728 VDD CLK 367 VDD P12LL L=6E-08 W=1E-06 $X=17715 $Y=-100 $D=2
M729 VDD 196 103 VDD P12LL L=6E-08 W=2.5E-06 $X=17745 $Y=6890 $D=2
M730 200 197 VDD VDD P12LL L=6E-08 W=1E-06 $X=17985 $Y=-100 $D=2
M731 98 199 VDD VDD P12LL L=6E-08 W=4E-07 $X=17985 $Y=24010 $D=2
M732 YX[3] 199 58 VDD P12LL L=6E-08 W=1.25E-06 $X=17985 $Y=27205 $D=2
M733 YX[3] 98 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=17985 $Y=30765 $D=2
M734 103 196 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=18015 $Y=6890 $D=2
M735 207 99 VDD VDD P12LL L=1.5E-07 W=7E-07 $X=18035 $Y=10600 $D=2
M736 211 226 VDD VDD P12LL L=6E-08 W=1E-06 $X=18145 $Y=16080 $D=2
M737 201 ACTRCLK 199 VDD P12LL L=6E-08 W=5E-07 $X=18145 $Y=22055 $D=2
M738 215 198 58 VDD P12LL L=6E-08 W=5E-07 $X=18180 $Y=33805 $D=2
M739 58 198 215 VDD P12LL L=6E-08 W=5E-07 $X=18180 $Y=34075 $D=2
M740 VDD 71 201 VDD P12LL L=6E-08 W=1E-06 $X=18275 $Y=17910 $D=2
M741 VDD 199 98 VDD P12LL L=6E-08 W=4E-07 $X=18275 $Y=24010 $D=2
M742 58 199 YX[3] VDD P12LL L=6E-08 W=1.25E-06 $X=18275 $Y=27205 $D=2
M743 VDD 98 YX[3] VDD P12LL L=6E-08 W=1.25E-06 $X=18275 $Y=30765 $D=2
M744 VDD 196 103 VDD P12LL L=6E-08 W=2.5E-06 $X=18285 $Y=6890 $D=2
M745 VDD 226 211 VDD P12LL L=6E-08 W=1E-06 $X=18415 $Y=16080 $D=2
M746 199 ACTRCLK 201 VDD P12LL L=6E-08 W=5E-07 $X=18415 $Y=22055 $D=2
M747 VDD 98 199 VDD P12LL L=3E-07 W=1.2E-07 $X=18525 $Y=23170 $D=2
M748 201 68 VDD VDD P12LL L=6E-08 W=1E-06 $X=18565 $Y=17910 $D=2
M749 98 199 VDD VDD P12LL L=6E-08 W=4E-07 $X=18565 $Y=24010 $D=2
M750 YX[3] 199 58 VDD P12LL L=6E-08 W=1.25E-06 $X=18565 $Y=27205 $D=2
M751 YX[3] 98 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=18565 $Y=30765 $D=2
M752 202 200 VDD VDD P12LL L=6E-08 W=1E-06 $X=18595 $Y=-100 $D=2
M753 201 ACTRCLK 199 VDD P12LL L=6E-08 W=5E-07 $X=18695 $Y=22055 $D=2
M754 226 205 VDD VDD P12LL L=6E-08 W=1E-06 $X=18705 $Y=16080 $D=2
M755 VDD 211 201 VDD P12LL L=6E-08 W=1E-06 $X=18855 $Y=17910 $D=2
M756 VDD 199 98 VDD P12LL L=6E-08 W=4E-07 $X=18855 $Y=24010 $D=2
M757 58 199 YX[3] VDD P12LL L=6E-08 W=1.25E-06 $X=18855 $Y=27205 $D=2
M758 VDD 98 YX[3] VDD P12LL L=6E-08 W=1.25E-06 $X=18855 $Y=30765 $D=2
M759 VDD 200 202 VDD P12LL L=6E-08 W=1E-06 $X=18865 $Y=-100 $D=2
M760 49 103 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=18895 $Y=6890 $D=2
M761 VDD 205 226 VDD P12LL L=6E-08 W=1E-06 $X=18995 $Y=16080 $D=2
M762 EMCLK 87 203 VDD P12LL L=6E-08 W=1.25E-06 $X=19115 $Y=10050 $D=2
M763 202 200 VDD VDD P12LL L=6E-08 W=1E-06 $X=19135 $Y=-100 $D=2
M764 102 211 VDD VDD P12LL L=6E-08 W=1E-06 $X=19145 $Y=17910 $D=2
M765 101 206 VDD VDD P12LL L=6E-08 W=4E-07 $X=19145 $Y=24010 $D=2
M766 YX[2] 206 58 VDD P12LL L=6E-08 W=1.25E-06 $X=19145 $Y=27205 $D=2
M767 YX[2] 101 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=19145 $Y=30765 $D=2
M768 VDD 103 49 VDD P12LL L=6E-08 W=2.5E-06 $X=19165 $Y=6890 $D=2
M769 215 209 VDD VDD P12LL L=6E-08 W=1E-06 $X=19180 $Y=33805 $D=2
M770 VDD 209 215 VDD P12LL L=6E-08 W=1E-06 $X=19180 $Y=34075 $D=2
M771 206 101 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=19235 $Y=23170 $D=2
M772 206 ACTRCLK 102 VDD P12LL L=6E-08 W=5E-07 $X=19305 $Y=22055 $D=2
M773 203 87 EMCLK VDD P12LL L=6E-08 W=1.25E-06 $X=19365 $Y=10050 $D=2
M774 49 103 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=19435 $Y=6890 $D=2
M775 VDD 68 102 VDD P12LL L=6E-08 W=1E-06 $X=19435 $Y=17910 $D=2
M776 VDD 206 101 VDD P12LL L=6E-08 W=4E-07 $X=19435 $Y=24010 $D=2
M777 58 206 YX[2] VDD P12LL L=6E-08 W=1.25E-06 $X=19435 $Y=27205 $D=2
M778 VDD 101 YX[2] VDD P12LL L=6E-08 W=1.25E-06 $X=19435 $Y=30765 $D=2
M779 102 ACTRCLK 206 VDD P12LL L=6E-08 W=5E-07 $X=19585 $Y=22055 $D=2
M780 368 YA[2] 205 VDD P12LL L=6E-08 W=4E-07 $X=19625 $Y=16410 $D=2
M781 VDD 103 49 VDD P12LL L=6E-08 W=2.5E-06 $X=19705 $Y=6890 $D=2
M782 VDD 207 203 VDD P12LL L=6E-08 W=1.4E-06 $X=19710 $Y=9900 $D=2
M783 102 67 VDD VDD P12LL L=6E-08 W=1E-06 $X=19725 $Y=17910 $D=2
M784 101 206 VDD VDD P12LL L=6E-08 W=4E-07 $X=19725 $Y=24010 $D=2
M785 YX[2] 206 58 VDD P12LL L=6E-08 W=1.25E-06 $X=19725 $Y=27205 $D=2
M786 YX[2] 101 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=19725 $Y=30765 $D=2
M787 206 ACTRCLK 102 VDD P12LL L=6E-08 W=5E-07 $X=19855 $Y=22055 $D=2
M788 VDD VSS 368 VDD P12LL L=1E-07 W=4E-07 $X=19915 $Y=16410 $D=2
M789 49 103 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=19975 $Y=6890 $D=2
M790 99 212 VDD VDD P12LL L=6E-08 W=1.4E-06 $X=19980 $Y=9900 $D=2
M791 VDD 206 101 VDD P12LL L=6E-08 W=4E-07 $X=20015 $Y=24010 $D=2
M792 58 206 YX[2] VDD P12LL L=6E-08 W=1.25E-06 $X=20015 $Y=27205 $D=2
M793 VDD 101 YX[2] VDD P12LL L=6E-08 W=1.25E-06 $X=20015 $Y=30765 $D=2
M794 VDD 49 103 VDD P12LL L=2E-07 W=1.2E-07 $X=20125 $Y=-105 $D=2
M795 VDD 213 220 VDD P12LL L=2E-07 W=4E-07 $X=20145 $Y=680 $D=2
M796 VDD 103 49 VDD P12LL L=6E-08 W=2.5E-06 $X=20245 $Y=6890 $D=2
M797 105 210 VDD VDD P12LL L=6E-08 W=4E-07 $X=20305 $Y=24010 $D=2
M798 YX[0] 210 58 VDD P12LL L=6E-08 W=1.25E-06 $X=20305 $Y=27205 $D=2
M799 YX[0] 105 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=20305 $Y=30765 $D=2
M800 EMCLK 83 99 VDD P12LL L=6E-08 W=1.25E-06 $X=20320 $Y=10050 $D=2
M801 104 ACTRCLK 210 VDD P12LL L=6E-08 W=5E-07 $X=20465 $Y=22055 $D=2
M802 49 103 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=20515 $Y=6890 $D=2
M803 99 83 EMCLK VDD P12LL L=6E-08 W=1.25E-06 $X=20570 $Y=10050 $D=2
M804 VDD 67 104 VDD P12LL L=6E-08 W=1E-06 $X=20595 $Y=17910 $D=2
M805 VDD 210 105 VDD P12LL L=6E-08 W=4E-07 $X=20595 $Y=24010 $D=2
M806 58 210 YX[0] VDD P12LL L=6E-08 W=1.25E-06 $X=20595 $Y=27205 $D=2
M807 VDD 105 YX[0] VDD P12LL L=6E-08 W=1.25E-06 $X=20595 $Y=30765 $D=2
M808 369 VSS VDD VDD P12LL L=2E-07 W=8E-07 $X=20615 $Y=380 $D=2
M809 210 ACTRCLK 104 VDD P12LL L=6E-08 W=5E-07 $X=20735 $Y=22055 $D=2
M810 VDD 103 49 VDD P12LL L=6E-08 W=2.5E-06 $X=20785 $Y=6890 $D=2
M811 VDD 105 210 VDD P12LL L=3E-07 W=1.2E-07 $X=20845 $Y=23170 $D=2
M812 104 230 VDD VDD P12LL L=6E-08 W=1E-06 $X=20885 $Y=17910 $D=2
M813 105 210 VDD VDD P12LL L=6E-08 W=4E-07 $X=20885 $Y=24010 $D=2
M814 YX[0] 210 58 VDD P12LL L=6E-08 W=1.25E-06 $X=20885 $Y=27205 $D=2
M815 YX[0] 105 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=20885 $Y=30765 $D=2
M816 104 ACTRCLK 210 VDD P12LL L=6E-08 W=5E-07 $X=21015 $Y=22055 $D=2
M817 213 49 369 VDD P12LL L=2E-07 W=8E-07 $X=21065 $Y=380 $D=2
M818 58 49 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=21075 $Y=6890 $D=2
M819 VDD 211 104 VDD P12LL L=6E-08 W=1E-06 $X=21175 $Y=17910 $D=2
M820 VDD 210 105 VDD P12LL L=6E-08 W=4E-07 $X=21175 $Y=24010 $D=2
M821 58 210 YX[0] VDD P12LL L=6E-08 W=1.25E-06 $X=21175 $Y=27205 $D=2
M822 VDD 105 YX[0] VDD P12LL L=6E-08 W=1.25E-06 $X=21175 $Y=30765 $D=2
M823 VDD 218 212 VDD P12LL L=1.5E-07 W=7E-07 $X=21315 $Y=10600 $D=2
M824 VDD 49 58 VDD P12LL L=6E-08 W=2.5E-06 $X=21345 $Y=6890 $D=2
M825 216 211 VDD VDD P12LL L=6E-08 W=1E-06 $X=21465 $Y=17910 $D=2
M826 106 214 VDD VDD P12LL L=6E-08 W=4E-07 $X=21465 $Y=24010 $D=2
M827 YX[1] 214 58 VDD P12LL L=6E-08 W=1.25E-06 $X=21465 $Y=27205 $D=2
M828 YX[1] 106 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=21465 $Y=30765 $D=2
M829 214 106 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=21555 $Y=23170 $D=2
M830 58 49 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=21615 $Y=6890 $D=2
M831 214 ACTRCLK 216 VDD P12LL L=6E-08 W=5E-07 $X=21625 $Y=22055 $D=2
M832 VDD 230 216 VDD P12LL L=6E-08 W=1E-06 $X=21755 $Y=17910 $D=2
M833 VDD 214 106 VDD P12LL L=6E-08 W=4E-07 $X=21755 $Y=24010 $D=2
M834 58 214 YX[1] VDD P12LL L=6E-08 W=1.25E-06 $X=21755 $Y=27205 $D=2
M835 VDD 106 YX[1] VDD P12LL L=6E-08 W=1.25E-06 $X=21755 $Y=30765 $D=2
M836 370 VSS VDD VDD P12LL L=1E-07 W=4E-07 $X=21825 $Y=16410 $D=2
M837 VDD 49 58 VDD P12LL L=6E-08 W=2.5E-06 $X=21885 $Y=6890 $D=2
M838 VDD 49 217 VDD P12LL L=2E-07 W=4E-07 $X=21895 $Y=680 $D=2
M839 216 ACTRCLK 214 VDD P12LL L=6E-08 W=5E-07 $X=21905 $Y=22055 $D=2
M840 216 71 VDD VDD P12LL L=6E-08 W=1E-06 $X=22045 $Y=17910 $D=2
M841 106 214 VDD VDD P12LL L=6E-08 W=4E-07 $X=22045 $Y=24010 $D=2
M842 YX[1] 214 58 VDD P12LL L=6E-08 W=1.25E-06 $X=22045 $Y=27205 $D=2
M843 YX[1] 106 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=22045 $Y=30765 $D=2
M844 EMCLK 183 218 VDD P12LL L=6E-08 W=1E-06 $X=22060 $Y=10400 $D=2
M845 219 YA[0] 370 VDD P12LL L=6E-08 W=4E-07 $X=22155 $Y=16410 $D=2
M846 214 ACTRCLK 216 VDD P12LL L=6E-08 W=5E-07 $X=22175 $Y=22055 $D=2
M847 218 183 EMCLK VDD P12LL L=6E-08 W=1E-06 $X=22330 $Y=10400 $D=2
M848 VDD 214 106 VDD P12LL L=6E-08 W=4E-07 $X=22335 $Y=24010 $D=2
M849 58 214 YX[1] VDD P12LL L=6E-08 W=1.25E-06 $X=22335 $Y=27205 $D=2
M850 VDD 106 YX[1] VDD P12LL L=6E-08 W=1.25E-06 $X=22335 $Y=30765 $D=2
M851 223 217 VDD VDD P12LL L=2E-07 W=4E-07 $X=22385 $Y=680 $D=2
M852 108 222 VDD VDD P12LL L=6E-08 W=4E-07 $X=22625 $Y=24010 $D=2
M853 YX[7] 222 58 VDD P12LL L=6E-08 W=1.25E-06 $X=22625 $Y=27205 $D=2
M854 YX[7] 108 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=22625 $Y=30765 $D=2
M855 VDD 221 218 VDD P12LL L=6E-08 W=1.4E-06 $X=22645 $Y=10000 $D=2
M856 71 219 VDD VDD P12LL L=6E-08 W=1E-06 $X=22785 $Y=16080 $D=2
M857 107 ACTRCLK 222 VDD P12LL L=6E-08 W=5E-07 $X=22785 $Y=22055 $D=2
M858 221 103 VDD VDD P12LL L=6E-08 W=1.4E-06 $X=22915 $Y=10000 $D=2
M859 VDD 71 107 VDD P12LL L=6E-08 W=1E-06 $X=22915 $Y=17910 $D=2
M860 VDD 222 108 VDD P12LL L=6E-08 W=4E-07 $X=22915 $Y=24010 $D=2
M861 58 222 YX[7] VDD P12LL L=6E-08 W=1.25E-06 $X=22915 $Y=27205 $D=2
M862 VDD 108 YX[7] VDD P12LL L=6E-08 W=1.25E-06 $X=22915 $Y=30765 $D=2
M863 222 ACTRCLK 107 VDD P12LL L=6E-08 W=5E-07 $X=23055 $Y=22055 $D=2
M864 VDD 219 71 VDD P12LL L=6E-08 W=1E-06 $X=23075 $Y=16080 $D=2
M865 371 49 109 VDD P12LL L=6E-08 W=1.5E-06 $X=23125 $Y=-365 $D=2
M866 VDD 108 222 VDD P12LL L=3E-07 W=1.2E-07 $X=23165 $Y=23170 $D=2
M867 107 68 VDD VDD P12LL L=6E-08 W=1E-06 $X=23205 $Y=17910 $D=2
M868 108 222 VDD VDD P12LL L=6E-08 W=4E-07 $X=23205 $Y=24010 $D=2
M869 YX[7] 222 58 VDD P12LL L=6E-08 W=1.25E-06 $X=23205 $Y=27205 $D=2
M870 YX[7] 108 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=23205 $Y=30765 $D=2
M871 107 ACTRCLK 222 VDD P12LL L=6E-08 W=5E-07 $X=23335 $Y=22055 $D=2
M872 67 71 VDD VDD P12LL L=6E-08 W=1E-06 $X=23365 $Y=16080 $D=2
M873 VDD 223 371 VDD P12LL L=6E-08 W=1.5E-06 $X=23395 $Y=-365 $D=2
M874 VDD 226 107 VDD P12LL L=6E-08 W=1E-06 $X=23495 $Y=17910 $D=2
M875 VDD 222 108 VDD P12LL L=6E-08 W=4E-07 $X=23495 $Y=24010 $D=2
M876 58 222 YX[7] VDD P12LL L=6E-08 W=1.25E-06 $X=23495 $Y=27205 $D=2
M877 VDD 108 YX[7] VDD P12LL L=6E-08 W=1.25E-06 $X=23495 $Y=30765 $D=2
M878 VDD 71 67 VDD P12LL L=6E-08 W=1E-06 $X=23635 $Y=16080 $D=2
M879 372 223 VDD VDD P12LL L=6E-08 W=1.5E-06 $X=23665 $Y=-365 $D=2
M880 110 226 VDD VDD P12LL L=6E-08 W=1E-06 $X=23785 $Y=17910 $D=2
M881 111 224 VDD VDD P12LL L=6E-08 W=4E-07 $X=23785 $Y=24010 $D=2
M882 YX[6] 224 58 VDD P12LL L=6E-08 W=1.25E-06 $X=23785 $Y=27205 $D=2
M883 YX[6] 111 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=23785 $Y=30765 $D=2
M884 RWLR 215 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=23810 $Y=33805 $D=2
M885 VDD 215 RWLR VDD P12LL L=6E-08 W=2.5E-06 $X=23810 $Y=34075 $D=2
M886 224 111 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=23875 $Y=23170 $D=2
M887 SACK1 49 VDD VDD P12LL L=6E-08 W=5E-06 $X=23925 $Y=4275 $D=2
M888 109 49 372 VDD P12LL L=6E-08 W=1.5E-06 $X=23935 $Y=-365 $D=2
M889 224 ACTRCLK 110 VDD P12LL L=6E-08 W=5E-07 $X=23945 $Y=22055 $D=2
M890 VDD 68 110 VDD P12LL L=6E-08 W=1E-06 $X=24075 $Y=17910 $D=2
M891 VDD 224 111 VDD P12LL L=6E-08 W=4E-07 $X=24075 $Y=24010 $D=2
M892 58 224 YX[6] VDD P12LL L=6E-08 W=1.25E-06 $X=24075 $Y=27205 $D=2
M893 VDD 111 YX[6] VDD P12LL L=6E-08 W=1.25E-06 $X=24075 $Y=30765 $D=2
M894 VDD 49 SACK1 VDD P12LL L=6E-08 W=5E-06 $X=24195 $Y=4275 $D=2
M895 110 ACTRCLK 224 VDD P12LL L=6E-08 W=5E-07 $X=24225 $Y=22055 $D=2
M896 110 67 VDD VDD P12LL L=6E-08 W=1E-06 $X=24365 $Y=17910 $D=2
M897 111 224 VDD VDD P12LL L=6E-08 W=4E-07 $X=24365 $Y=24010 $D=2
M898 YX[6] 224 58 VDD P12LL L=6E-08 W=1.25E-06 $X=24365 $Y=27205 $D=2
M899 YX[6] 111 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=24365 $Y=30765 $D=2
M900 SACK4 109 VDD VDD P12LL L=6E-08 W=5E-06 $X=24465 $Y=4275 $D=2
M901 224 ACTRCLK 110 VDD P12LL L=6E-08 W=5E-07 $X=24495 $Y=22055 $D=2
M902 373 220 228 VDD P12LL L=6E-08 W=1.25E-06 $X=24545 $Y=-115 $D=2
M903 VDD 224 111 VDD P12LL L=6E-08 W=4E-07 $X=24655 $Y=24010 $D=2
M904 58 224 YX[6] VDD P12LL L=6E-08 W=1.25E-06 $X=24655 $Y=27205 $D=2
M905 VDD 111 YX[6] VDD P12LL L=6E-08 W=1.25E-06 $X=24655 $Y=30765 $D=2
M906 VDD 109 SACK4 VDD P12LL L=6E-08 W=5E-06 $X=24735 $Y=4275 $D=2
M907 VDD 49 373 VDD P12LL L=6E-08 W=1.25E-06 $X=24815 $Y=-115 $D=2
M908 112 225 VDD VDD P12LL L=6E-08 W=4E-07 $X=24945 $Y=24010 $D=2
M909 YX[4] 225 58 VDD P12LL L=6E-08 W=1.25E-06 $X=24945 $Y=27205 $D=2
M910 YX[4] 112 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=24945 $Y=30765 $D=2
M911 DCTRCLK 228 VDD VDD P12LL L=6E-08 W=5E-06 $X=25005 $Y=4275 $D=2
M912 374 VSS VDD VDD P12LL L=1E-07 W=4E-07 $X=25005 $Y=16410 $D=2
M913 375 49 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=25085 $Y=-115 $D=2
M914 113 ACTRCLK 225 VDD P12LL L=6E-08 W=5E-07 $X=25105 $Y=22055 $D=2
M915 VDD 67 113 VDD P12LL L=6E-08 W=1E-06 $X=25235 $Y=17910 $D=2
M916 VDD 225 112 VDD P12LL L=6E-08 W=4E-07 $X=25235 $Y=24010 $D=2
M917 58 225 YX[4] VDD P12LL L=6E-08 W=1.25E-06 $X=25235 $Y=27205 $D=2
M918 VDD 112 YX[4] VDD P12LL L=6E-08 W=1.25E-06 $X=25235 $Y=30765 $D=2
M919 VDD 228 DCTRCLK VDD P12LL L=6E-08 W=5E-06 $X=25275 $Y=4275 $D=2
M920 227 YA[1] 374 VDD P12LL L=6E-08 W=4E-07 $X=25335 $Y=16410 $D=2
M921 228 220 375 VDD P12LL L=6E-08 W=1.25E-06 $X=25355 $Y=-115 $D=2
M922 225 ACTRCLK 113 VDD P12LL L=6E-08 W=5E-07 $X=25375 $Y=22055 $D=2
M923 VDD 112 225 VDD P12LL L=3E-07 W=1.2E-07 $X=25485 $Y=23170 $D=2
M924 113 230 VDD VDD P12LL L=6E-08 W=1E-06 $X=25525 $Y=17910 $D=2
M925 112 225 VDD VDD P12LL L=6E-08 W=4E-07 $X=25525 $Y=24010 $D=2
M926 YX[4] 225 58 VDD P12LL L=6E-08 W=1.25E-06 $X=25525 $Y=27205 $D=2
M927 YX[4] 112 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=25525 $Y=30765 $D=2
M928 ACTRCLK 228 VDD VDD P12LL L=6E-08 W=5E-06 $X=25545 $Y=4275 $D=2
M929 113 ACTRCLK 225 VDD P12LL L=6E-08 W=5E-07 $X=25655 $Y=22055 $D=2
M930 VDD 228 ACTRCLK VDD P12LL L=6E-08 W=5E-06 $X=25815 $Y=4275 $D=2
M931 VDD 226 113 VDD P12LL L=6E-08 W=1E-06 $X=25815 $Y=17910 $D=2
M932 VDD 225 112 VDD P12LL L=6E-08 W=4E-07 $X=25815 $Y=24010 $D=2
M933 58 225 YX[4] VDD P12LL L=6E-08 W=1.25E-06 $X=25815 $Y=27205 $D=2
M934 VDD 112 YX[4] VDD P12LL L=6E-08 W=1.25E-06 $X=25815 $Y=30765 $D=2
M935 231 228 VDD VDD P12LL L=6E-08 W=1E-06 $X=25945 $Y=70 $D=2
M936 68 227 VDD VDD P12LL L=6E-08 W=1E-06 $X=25965 $Y=16080 $D=2
M937 ACTRCLKX ACTRCLK VDD VDD P12LL L=6E-08 W=5E-06 $X=26085 $Y=4275 $D=2
M938 232 226 VDD VDD P12LL L=6E-08 W=1E-06 $X=26105 $Y=17910 $D=2
M939 114 229 VDD VDD P12LL L=6E-08 W=4E-07 $X=26105 $Y=24010 $D=2
M940 YX[5] 229 58 VDD P12LL L=6E-08 W=1.25E-06 $X=26105 $Y=27205 $D=2
M941 YX[5] 114 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=26105 $Y=30765 $D=2
M942 229 114 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=26195 $Y=23170 $D=2
M943 VDD 228 231 VDD P12LL L=6E-08 W=1E-06 $X=26215 $Y=70 $D=2
M944 VDD 227 68 VDD P12LL L=6E-08 W=1E-06 $X=26255 $Y=16080 $D=2
M945 229 ACTRCLK 232 VDD P12LL L=6E-08 W=5E-07 $X=26265 $Y=22055 $D=2
M946 VDD ACTRCLK ACTRCLKX VDD P12LL L=6E-08 W=5E-06 $X=26355 $Y=4275 $D=2
M947 VDD 230 232 VDD P12LL L=6E-08 W=1E-06 $X=26395 $Y=17910 $D=2
M948 VDD 229 114 VDD P12LL L=6E-08 W=4E-07 $X=26395 $Y=24010 $D=2
M949 58 229 YX[5] VDD P12LL L=6E-08 W=1.25E-06 $X=26395 $Y=27205 $D=2
M950 VDD 114 YX[5] VDD P12LL L=6E-08 W=1.25E-06 $X=26395 $Y=30765 $D=2
M951 231 228 VDD VDD P12LL L=6E-08 W=1E-06 $X=26485 $Y=70 $D=2
M952 230 68 VDD VDD P12LL L=6E-08 W=1E-06 $X=26545 $Y=16080 $D=2
M953 232 ACTRCLK 229 VDD P12LL L=6E-08 W=5E-07 $X=26545 $Y=22055 $D=2
M954 DCTRCLKX 231 VDD VDD P12LL L=6E-08 W=5E-06 $X=26625 $Y=4275 $D=2
M955 232 71 VDD VDD P12LL L=6E-08 W=1E-06 $X=26685 $Y=17910 $D=2
M956 114 229 VDD VDD P12LL L=6E-08 W=4E-07 $X=26685 $Y=24010 $D=2
M957 YX[5] 229 58 VDD P12LL L=6E-08 W=1.25E-06 $X=26685 $Y=27205 $D=2
M958 YX[5] 114 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=26685 $Y=30765 $D=2
M959 VDD 68 230 VDD P12LL L=6E-08 W=1E-06 $X=26815 $Y=16080 $D=2
M960 229 ACTRCLK 232 VDD P12LL L=6E-08 W=5E-07 $X=26815 $Y=22055 $D=2
M961 VDD 231 DCTRCLKX VDD P12LL L=6E-08 W=5E-06 $X=26895 $Y=4275 $D=2
M962 VDD 229 114 VDD P12LL L=6E-08 W=4E-07 $X=26975 $Y=24010 $D=2
M963 58 229 YX[5] VDD P12LL L=6E-08 W=1.25E-06 $X=26975 $Y=27205 $D=2
M964 VDD 114 YX[5] VDD P12LL L=6E-08 W=1.25E-06 $X=26975 $Y=30765 $D=2
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PYX
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PYX A CLK CLKX VDD VSS YAX
M0 38 36 VSS VSS N12LL L=6E-08 W=5E-07
M1 VSS 36 38 VSS N12LL L=6E-08 W=5E-07
M2 36 37 VSS VSS N12LL L=6E-08 W=4E-07
M3 1 CLKX 38 VSS N12LL L=6E-08 W=9E-07
M4 VSS 39 37 VSS N12LL L=3E-07 W=4E-07
M5 38 CLKX 1 VSS N12LL L=6E-08 W=8E-07
M6 39 A VSS VSS N12LL L=6E-08 W=4E-07
M7 1 CLKX 38 VSS N12LL L=6E-08 W=8E-07
M8 VSS YAX 1 VSS N12LL L=6E-07 W=1.2E-07
M9 YAX 1 VSS VSS N12LL L=6E-08 W=1E-06
M10 VSS 1 YAX VSS N12LL L=6E-08 W=1E-06
M11 YAX 1 VSS VSS N12LL L=6E-08 W=1E-06
M12 VSS 1 YAX VSS N12LL L=6E-08 W=1E-06
M13 YAX 1 VSS VSS N12LL L=6E-08 W=1E-06
M14 38 36 VDD VDD P12LL L=6E-08 W=1E-06
M15 VDD 36 38 VDD P12LL L=6E-08 W=1E-06
M16 36 37 VDD VDD P12LL L=6E-08 W=4E-07
M17 1 CLK 38 VDD P12LL L=6E-08 W=9E-07
M18 VDD 39 37 VDD P12LL L=3E-07 W=4E-07
M19 38 CLK 1 VDD P12LL L=6E-08 W=8E-07
M20 39 A VDD VDD P12LL L=6E-08 W=4E-07
M21 1 CLK 38 VDD P12LL L=6E-08 W=8E-07
M22 1 YAX VDD VDD P12LL L=3E-07 W=1.2E-07
M23 YAX 1 VDD VDD P12LL L=6E-08 W=2E-06
M24 VDD 1 YAX VDD P12LL L=6E-08 W=2E-06
M25 YAX 1 VDD VDD P12LL L=6E-08 W=2E-06
M26 VDD 1 YAX VDD P12LL L=6E-08 W=2E-06
M27 YAX 1 VDD VDD P12LL L=6E-08 W=2E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_LOGIC_BASEY16
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_LOGIC_BASEY16 ACTRCLK ACTRCLKX CEN CLK DCTRCLK DCTRCLKX EMCLK FB FCKX[7] FCKX[6]
+FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXA[2] PXA[1] PXA[0]
+RDE RWLL RWLR S[1] S[0] SACK1 SACK4 VDD VSS WE
+WEN XA[4] XA[3] XA[2] XA[1] XA[0] YA[3] YA[2] YA[1] YA[0]
+YAX YX[7] YX[6] YX[5] YX[4] YX[3] YX[2] YX[1] YX[0] ZA
+ZAX
XI0 RWLL RDE ACTRCLK ACTRCLKX ZAX PXA[3] PXA[2] PXA[1] PXA[0] XA[4]
+XA[3] XA[2] XA[1] XA[0] ZA FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3]
+FCKX[2] FCKX[1] FCKX[0] S[1] S[0] WEN WE CEN CLK FB
+YX[7] YX[6] YX[5] YX[4] YX[3] YX[2] YX[1] YX[0] YA[2] YA[1]
+YA[0] EMCLK RWLR SACK1 SACK4 DCTRCLK DCTRCLKX VDD VSS S55NLLGSPH_X512Y16D32_LOGIC_LEAFCELL_COMMON
XI1 YA[3] ACTRCLK ACTRCLKX VDD VSS YAX S55NLLGSPH_X512Y16D32_PYX
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_S65NLLHSDPH_ESDA12
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_S65NLLHSDPH_ESDA12 A[12] A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3]
+A[2] A[1] A[0] CEN CLK RDE S[1] S[0] VDD VSS
+WEN
MN12 A[12] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP12 VDD VDD A[12] VDD P12LL W=0.2U L=0.06U M=1
MN11 A[11] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP11 VDD VDD A[11] VDD P12LL W=0.2U L=0.06U M=1
MN10 A[10] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP10 VDD VDD A[10] VDD P12LL W=0.2U L=0.06U M=1
MN9 A[9] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP9 VDD VDD A[9] VDD P12LL W=0.2U L=0.06U M=1
MN8 A[8] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP8 VDD VDD A[8] VDD P12LL W=0.2U L=0.06U M=1
MN7 A[7] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP7 VDD VDD A[7] VDD P12LL W=0.2U L=0.06U M=1
MN6 A[6] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP6 VDD VDD A[6] VDD P12LL W=0.2U L=0.06U M=1
MN5 A[5] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP5 VDD VDD A[5] VDD P12LL W=0.2U L=0.06U M=1
MN4 A[4] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP4 VDD VDD A[4] VDD P12LL W=0.2U L=0.06U M=1
MN3 A[3] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP3 VDD VDD A[3] VDD P12LL W=0.2U L=0.06U M=1
MN2 A[2] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP2 VDD VDD A[2] VDD P12LL W=0.2U L=0.06U M=1
MN1 A[1] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP1 VDD VDD A[1] VDD P12LL W=0.2U L=0.06U M=1
MN0 A[0] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP0 VDD VDD A[0] VDD P12LL W=0.2U L=0.06U M=1
MN93 CEN VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MN91 WEN VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MN90 CLK VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP93 VDD VDD CEN VDD P12LL W=0.2U L=0.06U M=1
MP91 VDD VDD WEN VDD P12LL W=0.2U L=0.06U M=1
MP90 VDD VDD CLK VDD P12LL W=0.2U L=0.06U M=1
MM96 S[1] VSS VSS VSS N12LL W=200.0N L=60.00N M=1
MM98 S[0] VSS VSS VSS N12LL W=200.0N L=60.00N M=1
MM92 S[1] VDD VDD VDD P12LL W=200.0N L=60.00N M=1
MM94 S[0] VDD VDD VDD P12LL W=200.0N L=60.00N M=1
MM95 RDE VSS VSS VSS N12LL W=200.0N L=60.00N M=1
MM99 RDE VDD VDD VDD P12LL W=200.0N L=60.00N M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_TIE_LOW_X2
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_TIE_LOW_X2 VDD VSS PULL0
MN18 PULL0 NET18 VSS VSS N12LL W=1U L=60.00N M=1
MP18 NET18 NET18 VDD VDD P12LL W=400.0N L=60.00N M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_STWL_DEC
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_STWL_DEC EMCLK STWL VDD VSS
M0 2 5 VSS VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=1715 $D=0
M1 VSS 5 2 VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=1965 $D=0
M2 STWL 5 VSS VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=2215 $D=0
M3 VSS 5 STWL VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=2465 $D=0
M4 5 6 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=5800 $Y=2215 $D=0
M5 VSS 6 5 VSS N12LL L=6E-08 W=7.5E-07 $X=5800 $Y=2465 $D=0
M6 5 6 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=5800 $Y=2715 $D=0
M7 VSS 6 5 VSS N12LL L=6E-08 W=7.5E-07 $X=5800 $Y=2965 $D=0
M8 6 7 VSS VSS N12LL L=6E-08 W=8E-07 $X=9900 $Y=2220 $D=0
M9 7 12 EMCLK VSS N12LL L=6E-08 W=6E-07 $X=10020 $Y=2810 $D=0
M10 VSS 11 9 VSS N12LL L=6E-08 W=1E-06 $X=11775 $Y=2610 $D=0
M11 10 10 VSS VSS N12LL L=6E-08 W=4E-07 $X=12375 $Y=2930 $D=0
M12 2 5 VDD VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=1715 $D=14
M13 VDD 5 2 VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=1965 $D=14
M14 STWL 5 VDD VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=2215 $D=14
M15 VDD 5 STWL VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=2465 $D=14
M16 5 6 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=2215 $D=2
M17 VDD 6 5 VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=2465 $D=2
M18 5 6 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=2715 $D=2
M19 VDD 6 5 VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=2965 $D=2
M20 6 7 VDD VDD P12LL L=6E-08 W=4E-07 $X=8220 $Y=2220 $D=2
M21 VDD 7 6 VDD P12LL L=6E-08 W=4E-07 $X=8220 $Y=2485 $D=2
M22 7 9 EMCLK VDD P12LL L=6E-08 W=4E-07 $X=8960 $Y=2700 $D=2
M23 VDD 12 7 VDD P12LL L=6E-08 W=4E-07 $X=8960 $Y=2960 $D=2
M24 VDD 11 11 VDD P12LL L=6E-08 W=4E-07 $X=13570 $Y=2610 $D=2
M25 12 10 VDD VDD P12LL L=6E-08 W=1E-06 $X=13570 $Y=2930 $D=2
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_XDEC
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_XDEC FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA PXB
+PXC VDD VSS WLL[7] WLL[6] WLL[5] WLL[4] WLL[3] WLL[2] WLL[1]
+WLL[0] WLR[7] WLR[6] WLR[5] WLR[4] WLR[3] WLR[2] WLR[1] WLR[0]
M0 WLL[0] 11 VSS VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=695 $D=0
M1 VSS 11 WLL[0] VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=945 $D=0
M2 WLL[1] 12 VSS VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=1195 $D=0
M3 VSS 12 WLL[1] VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=1445 $D=0
M4 WLL[2] 13 VSS VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=1695 $D=0
M5 VSS 13 WLL[2] VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=1945 $D=0
M6 WLL[3] 14 VSS VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=2195 $D=0
M7 VSS 14 WLL[3] VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=2445 $D=0
M8 WLL[4] 15 VSS VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=2695 $D=0
M9 VSS 15 WLL[4] VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=2945 $D=0
M10 WLL[5] 16 VSS VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=3195 $D=0
M11 VSS 16 WLL[5] VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=3445 $D=0
M12 WLL[6] 17 VSS VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=3695 $D=0
M13 VSS 17 WLL[6] VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=3945 $D=0
M14 WLL[7] 18 VSS VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=4195 $D=0
M15 VSS 18 WLL[7] VSS N12LL L=6E-08 W=1E-06 $X=3890 $Y=4445 $D=0
M16 11 19 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=5780 $Y=695 $D=0
M17 VSS 19 11 VSS N12LL L=6E-08 W=7.5E-07 $X=5780 $Y=945 $D=0
M18 11 19 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=5780 $Y=1195 $D=0
M19 VSS 19 11 VSS N12LL L=6E-08 W=7.5E-07 $X=5780 $Y=1445 $D=0
M20 12 20 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=5780 $Y=1695 $D=0
M21 VSS 20 12 VSS N12LL L=6E-08 W=7.5E-07 $X=5780 $Y=1945 $D=0
M22 12 20 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=5780 $Y=2195 $D=0
M23 VSS 20 12 VSS N12LL L=6E-08 W=7.5E-07 $X=5780 $Y=2445 $D=0
M24 13 21 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=5780 $Y=2695 $D=0
M25 VSS 21 13 VSS N12LL L=6E-08 W=7.5E-07 $X=5780 $Y=2945 $D=0
M26 13 21 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=5780 $Y=3195 $D=0
M27 VSS 21 13 VSS N12LL L=6E-08 W=7.5E-07 $X=5780 $Y=3445 $D=0
M28 14 22 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=5780 $Y=3695 $D=0
M29 VSS 22 14 VSS N12LL L=6E-08 W=7.5E-07 $X=5780 $Y=3945 $D=0
M30 14 22 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=5780 $Y=4195 $D=0
M31 VSS 22 14 VSS N12LL L=6E-08 W=7.5E-07 $X=5780 $Y=4445 $D=0
M32 19 23 VSS VSS N12LL L=6E-08 W=8E-07 $X=9900 $Y=700 $D=0
M33 VSS 24 20 VSS N12LL L=6E-08 W=8E-07 $X=9900 $Y=2440 $D=0
M34 21 25 VSS VSS N12LL L=6E-08 W=8E-07 $X=9900 $Y=2700 $D=0
M35 VSS 26 22 VSS N12LL L=6E-08 W=8E-07 $X=9900 $Y=4440 $D=0
M36 23 35 FCKX[0] VSS N12LL L=6E-08 W=6E-07 $X=10020 $Y=1285 $D=0
M37 FCKX[1] 35 24 VSS N12LL L=6E-08 W=6E-07 $X=10020 $Y=1855 $D=0
M38 25 35 FCKX[2] VSS N12LL L=6E-08 W=6E-07 $X=10020 $Y=3285 $D=0
M39 FCKX[3] 35 26 VSS N12LL L=6E-08 W=6E-07 $X=10020 $Y=3855 $D=0
M40 36 35 VSS VSS N12LL L=6E-08 W=5E-07 $X=12815 $Y=1120 $D=0
M41 VSS 35 36 VSS N12LL L=6E-08 W=5E-07 $X=12815 $Y=1405 $D=0
M42 36 35 VSS VSS N12LL L=6E-08 W=5E-07 $X=12815 $Y=1695 $D=0
M43 VSS 35 36 VSS N12LL L=6E-08 W=5E-07 $X=12815 $Y=1985 $D=0
M44 35 34 VSS VSS N12LL L=6E-08 W=5E-07 $X=12815 $Y=2275 $D=0
M45 VSS 34 35 VSS N12LL L=6E-08 W=5E-07 $X=12815 $Y=2560 $D=0
M46 35 34 VSS VSS N12LL L=6E-08 W=5E-07 $X=12815 $Y=2850 $D=0
M47 VSS 34 35 VSS N12LL L=6E-08 W=5E-07 $X=12815 $Y=3140 $D=0
M48 88 PXA VSS VSS N12LL L=6E-08 W=8E-07 $X=12815 $Y=3430 $D=0
M49 89 PXB 88 VSS N12LL L=6E-08 W=8E-07 $X=12815 $Y=3720 $D=0
M50 34 PXC 89 VSS N12LL L=6E-08 W=8E-07 $X=12815 $Y=4010 $D=0
M51 45 41 VSS VSS N12LL L=6E-08 W=8E-07 $X=16550 $Y=700 $D=0
M52 VSS 42 46 VSS N12LL L=6E-08 W=8E-07 $X=16550 $Y=2440 $D=0
M53 47 43 VSS VSS N12LL L=6E-08 W=8E-07 $X=16550 $Y=2700 $D=0
M54 VSS 44 48 VSS N12LL L=6E-08 W=8E-07 $X=16550 $Y=4440 $D=0
M55 41 35 FCKX[4] VSS N12LL L=6E-08 W=6E-07 $X=16630 $Y=1290 $D=0
M56 FCKX[5] 35 42 VSS N12LL L=6E-08 W=6E-07 $X=16630 $Y=1850 $D=0
M57 43 35 FCKX[6] VSS N12LL L=6E-08 W=6E-07 $X=16630 $Y=3290 $D=0
M58 FCKX[7] 35 44 VSS N12LL L=6E-08 W=6E-07 $X=16630 $Y=3850 $D=0
M59 15 45 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=20720 $Y=695 $D=0
M60 VSS 45 15 VSS N12LL L=6E-08 W=7.5E-07 $X=20720 $Y=945 $D=0
M61 15 45 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=20720 $Y=1195 $D=0
M62 VSS 45 15 VSS N12LL L=6E-08 W=7.5E-07 $X=20720 $Y=1445 $D=0
M63 16 46 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=20720 $Y=1695 $D=0
M64 VSS 46 16 VSS N12LL L=6E-08 W=7.5E-07 $X=20720 $Y=1945 $D=0
M65 16 46 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=20720 $Y=2195 $D=0
M66 VSS 46 16 VSS N12LL L=6E-08 W=7.5E-07 $X=20720 $Y=2445 $D=0
M67 17 47 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=20720 $Y=2695 $D=0
M68 VSS 47 17 VSS N12LL L=6E-08 W=7.5E-07 $X=20720 $Y=2945 $D=0
M69 17 47 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=20720 $Y=3195 $D=0
M70 VSS 47 17 VSS N12LL L=6E-08 W=7.5E-07 $X=20720 $Y=3445 $D=0
M71 18 48 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=20720 $Y=3695 $D=0
M72 VSS 48 18 VSS N12LL L=6E-08 W=7.5E-07 $X=20720 $Y=3945 $D=0
M73 18 48 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=20720 $Y=4195 $D=0
M74 VSS 48 18 VSS N12LL L=6E-08 W=7.5E-07 $X=20720 $Y=4445 $D=0
M75 WLR[0] 11 VSS VSS N12LL L=6E-08 W=1E-06 $X=22360 $Y=695 $D=0
M76 VSS 11 WLR[0] VSS N12LL L=6E-08 W=1E-06 $X=22360 $Y=945 $D=0
M77 WLR[1] 12 VSS VSS N12LL L=6E-08 W=1E-06 $X=22360 $Y=1195 $D=0
M78 VSS 12 WLR[1] VSS N12LL L=6E-08 W=1E-06 $X=22360 $Y=1445 $D=0
M79 WLR[2] 13 VSS VSS N12LL L=6E-08 W=1E-06 $X=22360 $Y=1695 $D=0
M80 VSS 13 WLR[2] VSS N12LL L=6E-08 W=1E-06 $X=22360 $Y=1945 $D=0
M81 WLR[3] 14 VSS VSS N12LL L=6E-08 W=1E-06 $X=22360 $Y=2195 $D=0
M82 VSS 14 WLR[3] VSS N12LL L=6E-08 W=1E-06 $X=22360 $Y=2445 $D=0
M83 WLR[4] 15 VSS VSS N12LL L=6E-08 W=1E-06 $X=22360 $Y=2695 $D=0
M84 VSS 15 WLR[4] VSS N12LL L=6E-08 W=1E-06 $X=22360 $Y=2945 $D=0
M85 WLR[5] 16 VSS VSS N12LL L=6E-08 W=1E-06 $X=22360 $Y=3195 $D=0
M86 VSS 16 WLR[5] VSS N12LL L=6E-08 W=1E-06 $X=22360 $Y=3445 $D=0
M87 WLR[6] 17 VSS VSS N12LL L=6E-08 W=1E-06 $X=22360 $Y=3695 $D=0
M88 VSS 17 WLR[6] VSS N12LL L=6E-08 W=1E-06 $X=22360 $Y=3945 $D=0
M89 WLR[7] 18 VSS VSS N12LL L=6E-08 W=1E-06 $X=22360 $Y=4195 $D=0
M90 VSS 18 WLR[7] VSS N12LL L=6E-08 W=1E-06 $X=22360 $Y=4445 $D=0
M91 WLL[0] 11 VDD VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=695 $D=7
M92 VDD 11 WLL[0] VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=945 $D=7
M93 WLL[1] 12 VDD VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=1195 $D=7
M94 VDD 12 WLL[1] VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=1445 $D=7
M95 WLL[2] 13 VDD VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=1695 $D=7
M96 VDD 13 WLL[2] VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=1945 $D=7
M97 WLL[3] 14 VDD VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=2195 $D=7
M98 VDD 14 WLL[3] VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=2445 $D=7
M99 WLL[4] 15 VDD VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=2695 $D=7
M100 VDD 15 WLL[4] VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=2945 $D=7
M101 WLL[5] 16 VDD VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=3195 $D=7
M102 VDD 16 WLL[5] VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=3445 $D=7
M103 WLL[6] 17 VDD VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=3695 $D=7
M104 VDD 17 WLL[6] VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=3945 $D=7
M105 WLL[7] 18 VDD VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=4195 $D=7
M106 VDD 18 WLL[7] VDD PHVT12LL L=6E-08 W=2.5E-06 $X=940 $Y=4445 $D=7
M107 WLR[0] 11 VDD VDD PHVT12LL L=6E-08 W=2.5E-06 $X=23810 $Y=695 $D=7
M108 VDD 11 WLR[0] VDD PHVT12LL L=6E-08 W=2.5E-06 $X=23810 $Y=945 $D=7
M109 WLR[1] 12 VDD VDD PHVT12LL L=6E-08 W=2.5E-06 $X=23810 $Y=1195 $D=7
M110 VDD 12 WLR[1] VDD PHVT12LL L=6E-08 W=2.5E-06 $X=23810 $Y=1445 $D=7
M111 WLR[2] 13 VDD VDD PHVT12LL L=6E-08 W=2.5E-06 $X=23810 $Y=1695 $D=7
M112 VDD 13 WLR[2] VDD PHVT12LL L=6E-08 W=2.5E-06 $X=23810 $Y=1945 $D=7
M113 WLR[3] 14 VDD VDD PHVT12LL L=6E-08 W=2.5E-06 $X=23810 $Y=2195 $D=7
M114 VDD 14 WLR[3] VDD PHVT12LL L=6E-08 W=2.5E-06 $X=23810 $Y=2445 $D=7
M115 WLR[4] 15 VDD VDD PHVT12LL L=6E-08 W=2.5E-06 $X=23810 $Y=2695 $D=7
M116 VDD 15 WLR[4] VDD PHVT12LL L=6E-08 W=2.5E-06 $X=23810 $Y=2945 $D=7
M117 WLR[5] 16 VDD VDD PHVT12LL L=6E-08 W=2.5E-06 $X=23810 $Y=3195 $D=7
M118 VDD 16 WLR[5] VDD PHVT12LL L=6E-08 W=2.5E-06 $X=23810 $Y=3445 $D=7
M119 WLR[6] 17 VDD VDD PHVT12LL L=6E-08 W=2.5E-06 $X=23810 $Y=3695 $D=7
M120 VDD 17 WLR[6] VDD PHVT12LL L=6E-08 W=2.5E-06 $X=23810 $Y=3945 $D=7
M121 WLR[7] 18 VDD VDD PHVT12LL L=6E-08 W=2.5E-06 $X=23810 $Y=4195 $D=7
M122 VDD 18 WLR[7] VDD PHVT12LL L=6E-08 W=2.5E-06 $X=23810 $Y=4445 $D=7
M123 11 19 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=695 $D=1
M124 VDD 19 11 VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=945 $D=1
M125 11 19 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=1195 $D=1
M126 VDD 19 11 VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=1445 $D=1
M127 12 20 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=1695 $D=1
M128 VDD 20 12 VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=1945 $D=1
M129 12 20 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=2195 $D=1
M130 VDD 20 12 VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=2445 $D=1
M131 13 21 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=2695 $D=1
M132 VDD 21 13 VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=2945 $D=1
M133 13 21 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=3195 $D=1
M134 VDD 21 13 VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=3445 $D=1
M135 14 22 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=3695 $D=1
M136 VDD 22 14 VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=3945 $D=1
M137 14 22 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=4195 $D=1
M138 VDD 22 14 VDD P12LL L=6E-08 W=7.5E-07 $X=6950 $Y=4445 $D=1
M139 19 23 VDD VDD P12LL L=6E-08 W=4E-07 $X=8210 $Y=700 $D=1
M140 VDD 23 19 VDD P12LL L=6E-08 W=4E-07 $X=8210 $Y=965 $D=1
M141 20 24 VDD VDD P12LL L=6E-08 W=4E-07 $X=8210 $Y=2175 $D=1
M142 VDD 24 20 VDD P12LL L=6E-08 W=4E-07 $X=8210 $Y=2440 $D=1
M143 21 25 VDD VDD P12LL L=6E-08 W=4E-07 $X=8210 $Y=2700 $D=1
M144 VDD 25 21 VDD P12LL L=6E-08 W=4E-07 $X=8210 $Y=2965 $D=1
M145 22 26 VDD VDD P12LL L=6E-08 W=4E-07 $X=8210 $Y=4175 $D=1
M146 VDD 26 22 VDD P12LL L=6E-08 W=4E-07 $X=8210 $Y=4440 $D=1
M147 23 36 FCKX[0] VDD P12LL L=6E-08 W=4E-07 $X=8930 $Y=1180 $D=1
M148 VDD 35 23 VDD P12LL L=6E-08 W=4E-07 $X=8930 $Y=1440 $D=1
M149 24 35 VDD VDD P12LL L=6E-08 W=4E-07 $X=8930 $Y=1700 $D=1
M150 FCKX[1] 36 24 VDD P12LL L=6E-08 W=4E-07 $X=8930 $Y=1960 $D=1
M151 25 36 FCKX[2] VDD P12LL L=6E-08 W=4E-07 $X=8930 $Y=3180 $D=1
M152 VDD 35 25 VDD P12LL L=6E-08 W=4E-07 $X=8930 $Y=3440 $D=1
M153 26 35 VDD VDD P12LL L=6E-08 W=4E-07 $X=8930 $Y=3700 $D=1
M154 FCKX[3] 36 26 VDD P12LL L=6E-08 W=4E-07 $X=8930 $Y=3960 $D=1
M155 36 35 VDD VDD P12LL L=6E-08 W=5E-07 $X=14015 $Y=1120 $D=1
M156 VDD 35 36 VDD P12LL L=6E-08 W=5E-07 $X=14015 $Y=1405 $D=1
M157 36 35 VDD VDD P12LL L=6E-08 W=5E-07 $X=14015 $Y=1695 $D=1
M158 VDD 35 36 VDD P12LL L=6E-08 W=5E-07 $X=14015 $Y=1985 $D=1
M159 35 34 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=14015 $Y=2275 $D=1
M160 VDD 34 35 VDD P12LL L=6E-08 W=7.5E-07 $X=14015 $Y=2560 $D=1
M161 35 34 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=14015 $Y=2850 $D=1
M162 VDD 34 35 VDD P12LL L=6E-08 W=7.5E-07 $X=14015 $Y=3140 $D=1
M163 34 PXA VDD VDD P12LL L=6E-08 W=5E-07 $X=14015 $Y=3430 $D=1
M164 VDD PXB 34 VDD P12LL L=6E-08 W=5E-07 $X=14015 $Y=3720 $D=1
M165 34 PXC VDD VDD P12LL L=6E-08 W=5E-07 $X=14015 $Y=4010 $D=1
M166 41 36 FCKX[4] VDD P12LL L=6E-08 W=4E-07 $X=17920 $Y=1180 $D=1
M167 VDD 35 41 VDD P12LL L=6E-08 W=4E-07 $X=17920 $Y=1440 $D=1
M168 42 35 VDD VDD P12LL L=6E-08 W=4E-07 $X=17920 $Y=1700 $D=1
M169 FCKX[5] 36 42 VDD P12LL L=6E-08 W=4E-07 $X=17920 $Y=1960 $D=1
M170 43 36 FCKX[6] VDD P12LL L=6E-08 W=4E-07 $X=17920 $Y=3180 $D=1
M171 VDD 35 43 VDD P12LL L=6E-08 W=4E-07 $X=17920 $Y=3440 $D=1
M172 44 35 VDD VDD P12LL L=6E-08 W=4E-07 $X=17920 $Y=3700 $D=1
M173 FCKX[7] 36 44 VDD P12LL L=6E-08 W=4E-07 $X=17920 $Y=3960 $D=1
M174 45 41 VDD VDD P12LL L=6E-08 W=4E-07 $X=18640 $Y=700 $D=1
M175 VDD 41 45 VDD P12LL L=6E-08 W=4E-07 $X=18640 $Y=965 $D=1
M176 46 42 VDD VDD P12LL L=6E-08 W=4E-07 $X=18640 $Y=2175 $D=1
M177 VDD 42 46 VDD P12LL L=6E-08 W=4E-07 $X=18640 $Y=2440 $D=1
M178 47 43 VDD VDD P12LL L=6E-08 W=4E-07 $X=18640 $Y=2700 $D=1
M179 VDD 43 47 VDD P12LL L=6E-08 W=4E-07 $X=18640 $Y=2965 $D=1
M180 48 44 VDD VDD P12LL L=6E-08 W=4E-07 $X=18640 $Y=4175 $D=1
M181 VDD 44 48 VDD P12LL L=6E-08 W=4E-07 $X=18640 $Y=4440 $D=1
M182 15 45 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=19550 $Y=695 $D=1
M183 VDD 45 15 VDD P12LL L=6E-08 W=7.5E-07 $X=19550 $Y=945 $D=1
M184 15 45 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=19550 $Y=1195 $D=1
M185 VDD 45 15 VDD P12LL L=6E-08 W=7.5E-07 $X=19550 $Y=1445 $D=1
M186 16 46 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=19550 $Y=1695 $D=1
M187 VDD 46 16 VDD P12LL L=6E-08 W=7.5E-07 $X=19550 $Y=1945 $D=1
M188 16 46 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=19550 $Y=2195 $D=1
M189 VDD 46 16 VDD P12LL L=6E-08 W=7.5E-07 $X=19550 $Y=2445 $D=1
M190 17 47 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=19550 $Y=2695 $D=1
M191 VDD 47 17 VDD P12LL L=6E-08 W=7.5E-07 $X=19550 $Y=2945 $D=1
M192 17 47 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=19550 $Y=3195 $D=1
M193 VDD 47 17 VDD P12LL L=6E-08 W=7.5E-07 $X=19550 $Y=3445 $D=1
M194 18 48 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=19550 $Y=3695 $D=1
M195 VDD 48 18 VDD P12LL L=6E-08 W=7.5E-07 $X=19550 $Y=3945 $D=1
M196 18 48 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=19550 $Y=4195 $D=1
M197 VDD 48 18 VDD P12LL L=6E-08 W=7.5E-07 $X=19550 $Y=4445 $D=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_XDEC32
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_XDEC32 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXA[0]
+PXB[3] PXB[2] PXB[1] PXB[0] PXC[3] PXC[2] PXC[1] PXC[0] VDD VSS
+WLL[255] WLL[254] WLL[253] WLL[252] WLL[251] WLL[250] WLL[249] WLL[248] WLL[247] WLL[246]
+WLL[245] WLL[244] WLL[243] WLL[242] WLL[241] WLL[240] WLL[239] WLL[238] WLL[237] WLL[236]
+WLL[235] WLL[234] WLL[233] WLL[232] WLL[231] WLL[230] WLL[229] WLL[228] WLL[227] WLL[226]
+WLL[225] WLL[224] WLL[223] WLL[222] WLL[221] WLL[220] WLL[219] WLL[218] WLL[217] WLL[216]
+WLL[215] WLL[214] WLL[213] WLL[212] WLL[211] WLL[210] WLL[209] WLL[208] WLL[207] WLL[206]
+WLL[205] WLL[204] WLL[203] WLL[202] WLL[201] WLL[200] WLL[199] WLL[198] WLL[197] WLL[196]
+WLL[195] WLL[194] WLL[193] WLL[192] WLL[191] WLL[190] WLL[189] WLL[188] WLL[187] WLL[186]
+WLL[185] WLL[184] WLL[183] WLL[182] WLL[181] WLL[180] WLL[179] WLL[178] WLL[177] WLL[176]
+WLL[175] WLL[174] WLL[173] WLL[172] WLL[171] WLL[170] WLL[169] WLL[168] WLL[167] WLL[166]
+WLL[165] WLL[164] WLL[163] WLL[162] WLL[161] WLL[160] WLL[159] WLL[158] WLL[157] WLL[156]
+WLL[155] WLL[154] WLL[153] WLL[152] WLL[151] WLL[150] WLL[149] WLL[148] WLL[147] WLL[146]
+WLL[145] WLL[144] WLL[143] WLL[142] WLL[141] WLL[140] WLL[139] WLL[138] WLL[137] WLL[136]
+WLL[135] WLL[134] WLL[133] WLL[132] WLL[131] WLL[130] WLL[129] WLL[128] WLL[127] WLL[126]
+WLL[125] WLL[124] WLL[123] WLL[122] WLL[121] WLL[120] WLL[119] WLL[118] WLL[117] WLL[116]
+WLL[115] WLL[114] WLL[113] WLL[112] WLL[111] WLL[110] WLL[109] WLL[108] WLL[107] WLL[106]
+WLL[105] WLL[104] WLL[103] WLL[102] WLL[101] WLL[100] WLL[99] WLL[98] WLL[97] WLL[96]
+WLL[95] WLL[94] WLL[93] WLL[92] WLL[91] WLL[90] WLL[89] WLL[88] WLL[87] WLL[86]
+WLL[85] WLL[84] WLL[83] WLL[82] WLL[81] WLL[80] WLL[79] WLL[78] WLL[77] WLL[76]
+WLL[75] WLL[74] WLL[73] WLL[72] WLL[71] WLL[70] WLL[69] WLL[68] WLL[67] WLL[66]
+WLL[65] WLL[64] WLL[63] WLL[62] WLL[61] WLL[60] WLL[59] WLL[58] WLL[57] WLL[56]
+WLL[55] WLL[54] WLL[53] WLL[52] WLL[51] WLL[50] WLL[49] WLL[48] WLL[47] WLL[46]
+WLL[45] WLL[44] WLL[43] WLL[42] WLL[41] WLL[40] WLL[39] WLL[38] WLL[37] WLL[36]
+WLL[35] WLL[34] WLL[33] WLL[32] WLL[31] WLL[30] WLL[29] WLL[28] WLL[27] WLL[26]
+WLL[25] WLL[24] WLL[23] WLL[22] WLL[21] WLL[20] WLL[19] WLL[18] WLL[17] WLL[16]
+WLL[15] WLL[14] WLL[13] WLL[12] WLL[11] WLL[10] WLL[9] WLL[8] WLL[7] WLL[6]
+WLL[5] WLL[4] WLL[3] WLL[2] WLL[1] WLL[0] WLR[255] WLR[254] WLR[253] WLR[252]
+WLR[251] WLR[250] WLR[249] WLR[248] WLR[247] WLR[246] WLR[245] WLR[244] WLR[243] WLR[242]
+WLR[241] WLR[240] WLR[239] WLR[238] WLR[237] WLR[236] WLR[235] WLR[234] WLR[233] WLR[232]
+WLR[231] WLR[230] WLR[229] WLR[228] WLR[227] WLR[226] WLR[225] WLR[224] WLR[223] WLR[222]
+WLR[221] WLR[220] WLR[219] WLR[218] WLR[217] WLR[216] WLR[215] WLR[214] WLR[213] WLR[212]
+WLR[211] WLR[210] WLR[209] WLR[208] WLR[207] WLR[206] WLR[205] WLR[204] WLR[203] WLR[202]
+WLR[201] WLR[200] WLR[199] WLR[198] WLR[197] WLR[196] WLR[195] WLR[194] WLR[193] WLR[192]
+WLR[191] WLR[190] WLR[189] WLR[188] WLR[187] WLR[186] WLR[185] WLR[184] WLR[183] WLR[182]
+WLR[181] WLR[180] WLR[179] WLR[178] WLR[177] WLR[176] WLR[175] WLR[174] WLR[173] WLR[172]
+WLR[171] WLR[170] WLR[169] WLR[168] WLR[167] WLR[166] WLR[165] WLR[164] WLR[163] WLR[162]
+WLR[161] WLR[160] WLR[159] WLR[158] WLR[157] WLR[156] WLR[155] WLR[154] WLR[153] WLR[152]
+WLR[151] WLR[150] WLR[149] WLR[148] WLR[147] WLR[146] WLR[145] WLR[144] WLR[143] WLR[142]
+WLR[141] WLR[140] WLR[139] WLR[138] WLR[137] WLR[136] WLR[135] WLR[134] WLR[133] WLR[132]
+WLR[131] WLR[130] WLR[129] WLR[128] WLR[127] WLR[126] WLR[125] WLR[124] WLR[123] WLR[122]
+WLR[121] WLR[120] WLR[119] WLR[118] WLR[117] WLR[116] WLR[115] WLR[114] WLR[113] WLR[112]
+WLR[111] WLR[110] WLR[109] WLR[108] WLR[107] WLR[106] WLR[105] WLR[104] WLR[103] WLR[102]
+WLR[101] WLR[100] WLR[99] WLR[98] WLR[97] WLR[96] WLR[95] WLR[94] WLR[93] WLR[92]
+WLR[91] WLR[90] WLR[89] WLR[88] WLR[87] WLR[86] WLR[85] WLR[84] WLR[83] WLR[82]
+WLR[81] WLR[80] WLR[79] WLR[78] WLR[77] WLR[76] WLR[75] WLR[74] WLR[73] WLR[72]
+WLR[71] WLR[70] WLR[69] WLR[68] WLR[67] WLR[66] WLR[65] WLR[64] WLR[63] WLR[62]
+WLR[61] WLR[60] WLR[59] WLR[58] WLR[57] WLR[56] WLR[55] WLR[54] WLR[53] WLR[52]
+WLR[51] WLR[50] WLR[49] WLR[48] WLR[47] WLR[46] WLR[45] WLR[44] WLR[43] WLR[42]
+WLR[41] WLR[40] WLR[39] WLR[38] WLR[37] WLR[36] WLR[35] WLR[34] WLR[33] WLR[32]
+WLR[31] WLR[30] WLR[29] WLR[28] WLR[27] WLR[26] WLR[25] WLR[24] WLR[23] WLR[22]
+WLR[21] WLR[20] WLR[19] WLR[18] WLR[17] WLR[16] WLR[15] WLR[14] WLR[13] WLR[12]
+WLR[11] WLR[10] WLR[9] WLR[8] WLR[7] WLR[6] WLR[5] WLR[4] WLR[3] WLR[2]
+WLR[1] WLR[0]
XI0 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[3]
+PXC[3] VDD VSS WLL[255] WLL[254] WLL[253] WLL[252] WLL[251] WLL[250] WLL[249]
+WLL[248] WLR[255] WLR[254] WLR[253] WLR[252] WLR[251] WLR[250] WLR[249] WLR[248] S55NLLGSPH_X512Y16D32_XDEC
XI1 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[3]
+PXC[3] VDD VSS WLL[247] WLL[246] WLL[245] WLL[244] WLL[243] WLL[242] WLL[241]
+WLL[240] WLR[247] WLR[246] WLR[245] WLR[244] WLR[243] WLR[242] WLR[241] WLR[240] S55NLLGSPH_X512Y16D32_XDEC
XI2 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[2]
+PXC[3] VDD VSS WLL[239] WLL[238] WLL[237] WLL[236] WLL[235] WLL[234] WLL[233]
+WLL[232] WLR[239] WLR[238] WLR[237] WLR[236] WLR[235] WLR[234] WLR[233] WLR[232] S55NLLGSPH_X512Y16D32_XDEC
XI3 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[2]
+PXC[3] VDD VSS WLL[231] WLL[230] WLL[229] WLL[228] WLL[227] WLL[226] WLL[225]
+WLL[224] WLR[231] WLR[230] WLR[229] WLR[228] WLR[227] WLR[226] WLR[225] WLR[224] S55NLLGSPH_X512Y16D32_XDEC
XI4 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[1]
+PXC[3] VDD VSS WLL[223] WLL[222] WLL[221] WLL[220] WLL[219] WLL[218] WLL[217]
+WLL[216] WLR[223] WLR[222] WLR[221] WLR[220] WLR[219] WLR[218] WLR[217] WLR[216] S55NLLGSPH_X512Y16D32_XDEC
XI5 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[1]
+PXC[3] VDD VSS WLL[215] WLL[214] WLL[213] WLL[212] WLL[211] WLL[210] WLL[209]
+WLL[208] WLR[215] WLR[214] WLR[213] WLR[212] WLR[211] WLR[210] WLR[209] WLR[208] S55NLLGSPH_X512Y16D32_XDEC
XI6 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[0]
+PXC[3] VDD VSS WLL[207] WLL[206] WLL[205] WLL[204] WLL[203] WLL[202] WLL[201]
+WLL[200] WLR[207] WLR[206] WLR[205] WLR[204] WLR[203] WLR[202] WLR[201] WLR[200] S55NLLGSPH_X512Y16D32_XDEC
XI7 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[0]
+PXC[3] VDD VSS WLL[199] WLL[198] WLL[197] WLL[196] WLL[195] WLL[194] WLL[193]
+WLL[192] WLR[199] WLR[198] WLR[197] WLR[196] WLR[195] WLR[194] WLR[193] WLR[192] S55NLLGSPH_X512Y16D32_XDEC
XI8 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[3]
+PXC[2] VDD VSS WLL[191] WLL[190] WLL[189] WLL[188] WLL[187] WLL[186] WLL[185]
+WLL[184] WLR[191] WLR[190] WLR[189] WLR[188] WLR[187] WLR[186] WLR[185] WLR[184] S55NLLGSPH_X512Y16D32_XDEC
XI9 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[3]
+PXC[2] VDD VSS WLL[183] WLL[182] WLL[181] WLL[180] WLL[179] WLL[178] WLL[177]
+WLL[176] WLR[183] WLR[182] WLR[181] WLR[180] WLR[179] WLR[178] WLR[177] WLR[176] S55NLLGSPH_X512Y16D32_XDEC
XI10 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[2]
+PXC[2] VDD VSS WLL[175] WLL[174] WLL[173] WLL[172] WLL[171] WLL[170] WLL[169]
+WLL[168] WLR[175] WLR[174] WLR[173] WLR[172] WLR[171] WLR[170] WLR[169] WLR[168] S55NLLGSPH_X512Y16D32_XDEC
XI11 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[2]
+PXC[2] VDD VSS WLL[167] WLL[166] WLL[165] WLL[164] WLL[163] WLL[162] WLL[161]
+WLL[160] WLR[167] WLR[166] WLR[165] WLR[164] WLR[163] WLR[162] WLR[161] WLR[160] S55NLLGSPH_X512Y16D32_XDEC
XI12 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[1]
+PXC[2] VDD VSS WLL[159] WLL[158] WLL[157] WLL[156] WLL[155] WLL[154] WLL[153]
+WLL[152] WLR[159] WLR[158] WLR[157] WLR[156] WLR[155] WLR[154] WLR[153] WLR[152] S55NLLGSPH_X512Y16D32_XDEC
XI13 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[1]
+PXC[2] VDD VSS WLL[151] WLL[150] WLL[149] WLL[148] WLL[147] WLL[146] WLL[145]
+WLL[144] WLR[151] WLR[150] WLR[149] WLR[148] WLR[147] WLR[146] WLR[145] WLR[144] S55NLLGSPH_X512Y16D32_XDEC
XI14 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[0]
+PXC[2] VDD VSS WLL[143] WLL[142] WLL[141] WLL[140] WLL[139] WLL[138] WLL[137]
+WLL[136] WLR[143] WLR[142] WLR[141] WLR[140] WLR[139] WLR[138] WLR[137] WLR[136] S55NLLGSPH_X512Y16D32_XDEC
XI15 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[0]
+PXC[2] VDD VSS WLL[135] WLL[134] WLL[133] WLL[132] WLL[131] WLL[130] WLL[129]
+WLL[128] WLR[135] WLR[134] WLR[133] WLR[132] WLR[131] WLR[130] WLR[129] WLR[128] S55NLLGSPH_X512Y16D32_XDEC
XI16 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[3]
+PXC[1] VDD VSS WLL[127] WLL[126] WLL[125] WLL[124] WLL[123] WLL[122] WLL[121]
+WLL[120] WLR[127] WLR[126] WLR[125] WLR[124] WLR[123] WLR[122] WLR[121] WLR[120] S55NLLGSPH_X512Y16D32_XDEC
XI17 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[3]
+PXC[1] VDD VSS WLL[119] WLL[118] WLL[117] WLL[116] WLL[115] WLL[114] WLL[113]
+WLL[112] WLR[119] WLR[118] WLR[117] WLR[116] WLR[115] WLR[114] WLR[113] WLR[112] S55NLLGSPH_X512Y16D32_XDEC
XI18 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[2]
+PXC[1] VDD VSS WLL[111] WLL[110] WLL[109] WLL[108] WLL[107] WLL[106] WLL[105]
+WLL[104] WLR[111] WLR[110] WLR[109] WLR[108] WLR[107] WLR[106] WLR[105] WLR[104] S55NLLGSPH_X512Y16D32_XDEC
XI19 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[2]
+PXC[1] VDD VSS WLL[103] WLL[102] WLL[101] WLL[100] WLL[99] WLL[98] WLL[97]
+WLL[96] WLR[103] WLR[102] WLR[101] WLR[100] WLR[99] WLR[98] WLR[97] WLR[96] S55NLLGSPH_X512Y16D32_XDEC
XI20 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[1]
+PXC[1] VDD VSS WLL[95] WLL[94] WLL[93] WLL[92] WLL[91] WLL[90] WLL[89]
+WLL[88] WLR[95] WLR[94] WLR[93] WLR[92] WLR[91] WLR[90] WLR[89] WLR[88] S55NLLGSPH_X512Y16D32_XDEC
XI21 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[1]
+PXC[1] VDD VSS WLL[87] WLL[86] WLL[85] WLL[84] WLL[83] WLL[82] WLL[81]
+WLL[80] WLR[87] WLR[86] WLR[85] WLR[84] WLR[83] WLR[82] WLR[81] WLR[80] S55NLLGSPH_X512Y16D32_XDEC
XI22 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[0]
+PXC[1] VDD VSS WLL[79] WLL[78] WLL[77] WLL[76] WLL[75] WLL[74] WLL[73]
+WLL[72] WLR[79] WLR[78] WLR[77] WLR[76] WLR[75] WLR[74] WLR[73] WLR[72] S55NLLGSPH_X512Y16D32_XDEC
XI23 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[0]
+PXC[1] VDD VSS WLL[71] WLL[70] WLL[69] WLL[68] WLL[67] WLL[66] WLL[65]
+WLL[64] WLR[71] WLR[70] WLR[69] WLR[68] WLR[67] WLR[66] WLR[65] WLR[64] S55NLLGSPH_X512Y16D32_XDEC
XI24 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[3]
+PXC[0] VDD VSS WLL[63] WLL[62] WLL[61] WLL[60] WLL[59] WLL[58] WLL[57]
+WLL[56] WLR[63] WLR[62] WLR[61] WLR[60] WLR[59] WLR[58] WLR[57] WLR[56] S55NLLGSPH_X512Y16D32_XDEC
XI25 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[3]
+PXC[0] VDD VSS WLL[55] WLL[54] WLL[53] WLL[52] WLL[51] WLL[50] WLL[49]
+WLL[48] WLR[55] WLR[54] WLR[53] WLR[52] WLR[51] WLR[50] WLR[49] WLR[48] S55NLLGSPH_X512Y16D32_XDEC
XI26 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[2]
+PXC[0] VDD VSS WLL[47] WLL[46] WLL[45] WLL[44] WLL[43] WLL[42] WLL[41]
+WLL[40] WLR[47] WLR[46] WLR[45] WLR[44] WLR[43] WLR[42] WLR[41] WLR[40] S55NLLGSPH_X512Y16D32_XDEC
XI27 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[2]
+PXC[0] VDD VSS WLL[39] WLL[38] WLL[37] WLL[36] WLL[35] WLL[34] WLL[33]
+WLL[32] WLR[39] WLR[38] WLR[37] WLR[36] WLR[35] WLR[34] WLR[33] WLR[32] S55NLLGSPH_X512Y16D32_XDEC
XI28 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[1]
+PXC[0] VDD VSS WLL[31] WLL[30] WLL[29] WLL[28] WLL[27] WLL[26] WLL[25]
+WLL[24] WLR[31] WLR[30] WLR[29] WLR[28] WLR[27] WLR[26] WLR[25] WLR[24] S55NLLGSPH_X512Y16D32_XDEC
XI29 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[1]
+PXC[0] VDD VSS WLL[23] WLL[22] WLL[21] WLL[20] WLL[19] WLL[18] WLL[17]
+WLL[16] WLR[23] WLR[22] WLR[21] WLR[20] WLR[19] WLR[18] WLR[17] WLR[16] S55NLLGSPH_X512Y16D32_XDEC
XI30 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[0]
+PXC[0] VDD VSS WLL[15] WLL[14] WLL[13] WLL[12] WLL[11] WLL[10] WLL[9]
+WLL[8] WLR[15] WLR[14] WLR[13] WLR[12] WLR[11] WLR[10] WLR[9] WLR[8] S55NLLGSPH_X512Y16D32_XDEC
XI31 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[0]
+PXC[0] VDD VSS WLL[7] WLL[6] WLL[5] WLL[4] WLL[3] WLL[2] WLL[1]
+WLL[0] WLR[7] WLR[6] WLR[5] WLR[4] WLR[3] WLR[2] WLR[1] WLR[0] S55NLLGSPH_X512Y16D32_XDEC
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32_PX4
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32_PX4 A[0] A[1] CLK CLKX PX[3] PX[2] PX[1] PX[0] VDD VSS
M0 PX[3] 7 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=405 $Y=6825 $D=0
M1 12 PX[2] VSS VSS N12LL L=6E-07 W=1.2E-07 $X=485 $Y=6040 $D=0
M2 33 23 4 VSS N12LL L=6E-08 W=1.495E-06 $X=525 $Y=-4965 $D=0
M3 34 A[0] 5 VSS N12LL L=6E-08 W=4E-07 $X=545 $Y=-10675 $D=0
M4 7 CLKX 4 VSS N12LL L=6E-08 W=2.5E-06 $X=550 $Y=-725 $D=0
M5 VSS PX[3] 7 VSS N12LL L=6E-07 W=1.2E-07 $X=655 $Y=5355 $D=0
M6 VSS 7 PX[3] VSS N12LL L=6E-08 W=1.5E-06 $X=695 $Y=6825 $D=0
M7 VSS 17 33 VSS N12LL L=6E-08 W=1.495E-06 $X=705 $Y=-4965 $D=0
M8 VSS 5 23 VSS N12LL L=6E-08 W=7E-07 $X=740 $Y=-6515 $D=0
M9 VSS VDD 34 VSS N12LL L=3E-07 W=4E-07 $X=805 $Y=-10675 $D=0
M10 35 17 VSS VSS N12LL L=6E-08 W=1.495E-06 $X=975 $Y=-4965 $D=0
M11 PX[2] 12 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=985 $Y=6825 $D=0
M12 13 23 VSS VSS N12LL L=6E-08 W=7E-07 $X=1030 $Y=-6515 $D=0
M13 9 CLKX 12 VSS N12LL L=6E-08 W=2.5E-06 $X=1130 $Y=-725 $D=0
M14 9 13 35 VSS N12LL L=6E-08 W=1.495E-06 $X=1155 $Y=-4965 $D=0
M15 VSS 12 PX[2] VSS N12LL L=6E-08 W=1.5E-06 $X=1275 $Y=6825 $D=0
M16 PX[0] 14 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=1615 $Y=6825 $D=0
M17 21 PX[1] VSS VSS N12LL L=6E-07 W=1.2E-07 $X=1695 $Y=5355 $D=0
M18 36 13 15 VSS N12LL L=6E-08 W=1.495E-06 $X=1735 $Y=-4965 $D=0
M19 14 CLKX 15 VSS N12LL L=6E-08 W=2.5E-06 $X=1760 $Y=-725 $D=0
M20 VSS 22 17 VSS N12LL L=6E-08 W=7E-07 $X=1860 $Y=-6515 $D=0
M21 37 VDD VSS VSS N12LL L=3E-07 W=4E-07 $X=1865 $Y=-10675 $D=0
M22 VSS PX[0] 14 VSS N12LL L=6E-07 W=1.2E-07 $X=1865 $Y=6040 $D=0
M23 VSS 14 PX[0] VSS N12LL L=6E-08 W=1.5E-06 $X=1905 $Y=6825 $D=0
M24 VSS 20 36 VSS N12LL L=6E-08 W=1.495E-06 $X=1915 $Y=-4965 $D=0
M25 20 17 VSS VSS N12LL L=6E-08 W=7E-07 $X=2150 $Y=-6515 $D=0
M26 38 20 VSS VSS N12LL L=6E-08 W=1.495E-06 $X=2185 $Y=-4965 $D=0
M27 PX[1] 21 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=2195 $Y=6825 $D=0
M28 24 CLKX 21 VSS N12LL L=6E-08 W=2.5E-06 $X=2340 $Y=-725 $D=0
M29 22 A[1] 37 VSS N12LL L=6E-08 W=4E-07 $X=2365 $Y=-10675 $D=0
M30 24 23 38 VSS N12LL L=6E-08 W=1.495E-06 $X=2365 $Y=-4965 $D=0
M31 VSS 21 PX[1] VSS N12LL L=6E-08 W=1.5E-06 $X=2485 $Y=6825 $D=0
M32 PX[3] 7 VDD VDD P12LL L=6E-08 W=3.5E-06 $X=405 $Y=8930 $D=1
M33 4 23 VDD VDD P12LL L=6E-08 W=1.5E-06 $X=425 $Y=-2745 $D=1
M34 39 A[0] 5 VDD P12LL L=6E-08 W=4E-07 $X=545 $Y=-9440 $D=1
M35 7 CLK 4 VDD P12LL L=6E-08 W=2.5E-06 $X=550 $Y=2290 $D=1
M36 12 PX[2] VDD VDD P12LL L=3E-07 W=1.2E-07 $X=685 $Y=13080 $D=1
M37 VDD 7 PX[3] VDD P12LL L=6E-08 W=3.5E-06 $X=695 $Y=8930 $D=1
M38 VDD 17 4 VDD P12LL L=6E-08 W=1.5E-06 $X=705 $Y=-2745 $D=1
M39 VDD 5 23 VDD P12LL L=6E-08 W=1.4E-06 $X=740 $Y=-8525 $D=1
M40 VDD VSS 39 VDD P12LL L=1E-07 W=4E-07 $X=805 $Y=-9440 $D=1
M41 VDD PX[3] 7 VDD P12LL L=3E-07 W=1.2E-07 $X=940 $Y=13685 $D=1
M42 9 17 VDD VDD P12LL L=6E-08 W=1.5E-06 $X=975 $Y=-2745 $D=1
M43 PX[2] 12 VDD VDD P12LL L=6E-08 W=3.5E-06 $X=985 $Y=8930 $D=1
M44 13 23 VDD VDD P12LL L=6E-08 W=1.4E-06 $X=1030 $Y=-8525 $D=1
M45 9 CLK 12 VDD P12LL L=6E-08 W=2.5E-06 $X=1130 $Y=2290 $D=1
M46 VDD 13 9 VDD P12LL L=6E-08 W=1.5E-06 $X=1255 $Y=-2745 $D=1
M47 VDD 12 PX[2] VDD P12LL L=6E-08 W=3.5E-06 $X=1275 $Y=8930 $D=1
M48 PX[0] 14 VDD VDD P12LL L=6E-08 W=3.5E-06 $X=1615 $Y=8930 $D=1
M49 15 13 VDD VDD P12LL L=6E-08 W=1.5E-06 $X=1635 $Y=-2745 $D=1
M50 21 PX[1] VDD VDD P12LL L=3E-07 W=1.2E-07 $X=1710 $Y=13685 $D=1
M51 14 CLK 15 VDD P12LL L=6E-08 W=2.5E-06 $X=1760 $Y=2290 $D=1
M52 VDD 22 17 VDD P12LL L=6E-08 W=1.4E-06 $X=1860 $Y=-8525 $D=1
M53 VDD 14 PX[0] VDD P12LL L=6E-08 W=3.5E-06 $X=1905 $Y=8930 $D=1
M54 VDD 20 15 VDD P12LL L=6E-08 W=1.5E-06 $X=1915 $Y=-2745 $D=1
M55 VDD PX[0] 14 VDD P12LL L=3E-07 W=1.2E-07 $X=1965 $Y=13080 $D=1
M56 40 VSS VDD VDD P12LL L=1E-07 W=4E-07 $X=2065 $Y=-9440 $D=1
M57 20 17 VDD VDD P12LL L=6E-08 W=1.4E-06 $X=2150 $Y=-8525 $D=1
M58 24 20 VDD VDD P12LL L=6E-08 W=1.5E-06 $X=2185 $Y=-2745 $D=1
M59 PX[1] 21 VDD VDD P12LL L=6E-08 W=3.5E-06 $X=2195 $Y=8930 $D=1
M60 24 CLK 21 VDD P12LL L=6E-08 W=2.5E-06 $X=2340 $Y=2290 $D=1
M61 22 A[1] 40 VDD P12LL L=6E-08 W=4E-07 $X=2365 $Y=-9440 $D=1
M62 VDD 23 24 VDD P12LL L=6E-08 W=1.5E-06 $X=2465 $Y=-2745 $D=1
M63 VDD 21 PX[1] VDD P12LL L=6E-08 W=3.5E-06 $X=2485 $Y=8930 $D=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGSPH_X512Y16D32
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGSPH_X512Y16D32 A[12] A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3]
+A[2] A[1] A[0] CEN CLK D[31] D[30] D[29] D[28] D[27]
+D[26] D[25] D[24] D[23] D[22] D[21] D[20] D[19] D[18] D[17]
+D[16] D[15] D[14] D[13] D[12] D[11] D[10] D[9] D[8] D[7]
+D[6] D[5] D[4] D[3] D[2] D[1] D[0] Q[31] Q[30] Q[29]
+Q[28] Q[27] Q[26] Q[25] Q[24] Q[23] Q[22] Q[21] Q[20] Q[19]
+Q[18] Q[17] Q[16] Q[15] Q[14] Q[13] Q[12] Q[11] Q[10] Q[9]
+Q[8] Q[7] Q[6] Q[5] Q[4] Q[3] Q[2] Q[1] Q[0] VDD
+VSS WEN
XI0 D[15] D[14] D[13] D[12] D[11] D[10] D[9] D[8] D[7] D[6]
+D[5] D[4] D[3] D[2] D[1] D[0] DCTRCLK DCTRCLKX Q[15] Q[14]
+Q[13] Q[12] Q[11] Q[10] Q[9] Q[8] Q[7] Q[6] Q[5] Q[4]
+Q[3] Q[2] Q[1] Q[0] VSS VSS RWLL VSS SACK1 SACK4
+VSS VDD VSS WE WLL[511] WLL[510] WLL[509] WLL[508] WLL[507] WLL[506]
+WLL[505] WLL[504] WLL[503] WLL[502] WLL[501] WLL[500] WLL[499] WLL[498] WLL[497] WLL[496]
+WLL[495] WLL[494] WLL[493] WLL[492] WLL[491] WLL[490] WLL[489] WLL[488] WLL[487] WLL[486]
+WLL[485] WLL[484] WLL[483] WLL[482] WLL[481] WLL[480] WLL[479] WLL[478] WLL[477] WLL[476]
+WLL[475] WLL[474] WLL[473] WLL[472] WLL[471] WLL[470] WLL[469] WLL[468] WLL[467] WLL[466]
+WLL[465] WLL[464] WLL[463] WLL[462] WLL[461] WLL[460] WLL[459] WLL[458] WLL[457] WLL[456]
+WLL[455] WLL[454] WLL[453] WLL[452] WLL[451] WLL[450] WLL[449] WLL[448] WLL[447] WLL[446]
+WLL[445] WLL[444] WLL[443] WLL[442] WLL[441] WLL[440] WLL[439] WLL[438] WLL[437] WLL[436]
+WLL[435] WLL[434] WLL[433] WLL[432] WLL[431] WLL[430] WLL[429] WLL[428] WLL[427] WLL[426]
+WLL[425] WLL[424] WLL[423] WLL[422] WLL[421] WLL[420] WLL[419] WLL[418] WLL[417] WLL[416]
+WLL[415] WLL[414] WLL[413] WLL[412] WLL[411] WLL[410] WLL[409] WLL[408] WLL[407] WLL[406]
+WLL[405] WLL[404] WLL[403] WLL[402] WLL[401] WLL[400] WLL[399] WLL[398] WLL[397] WLL[396]
+WLL[395] WLL[394] WLL[393] WLL[392] WLL[391] WLL[390] WLL[389] WLL[388] WLL[387] WLL[386]
+WLL[385] WLL[384] WLL[383] WLL[382] WLL[381] WLL[380] WLL[379] WLL[378] WLL[377] WLL[376]
+WLL[375] WLL[374] WLL[373] WLL[372] WLL[371] WLL[370] WLL[369] WLL[368] WLL[367] WLL[366]
+WLL[365] WLL[364] WLL[363] WLL[362] WLL[361] WLL[360] WLL[359] WLL[358] WLL[357] WLL[356]
+WLL[355] WLL[354] WLL[353] WLL[352] WLL[351] WLL[350] WLL[349] WLL[348] WLL[347] WLL[346]
+WLL[345] WLL[344] WLL[343] WLL[342] WLL[341] WLL[340] WLL[339] WLL[338] WLL[337] WLL[336]
+WLL[335] WLL[334] WLL[333] WLL[332] WLL[331] WLL[330] WLL[329] WLL[328] WLL[327] WLL[326]
+WLL[325] WLL[324] WLL[323] WLL[322] WLL[321] WLL[320] WLL[319] WLL[318] WLL[317] WLL[316]
+WLL[315] WLL[314] WLL[313] WLL[312] WLL[311] WLL[310] WLL[309] WLL[308] WLL[307] WLL[306]
+WLL[305] WLL[304] WLL[303] WLL[302] WLL[301] WLL[300] WLL[299] WLL[298] WLL[297] WLL[296]
+WLL[295] WLL[294] WLL[293] WLL[292] WLL[291] WLL[290] WLL[289] WLL[288] WLL[287] WLL[286]
+WLL[285] WLL[284] WLL[283] WLL[282] WLL[281] WLL[280] WLL[279] WLL[278] WLL[277] WLL[276]
+WLL[275] WLL[274] WLL[273] WLL[272] WLL[271] WLL[270] WLL[269] WLL[268] WLL[267] WLL[266]
+WLL[265] WLL[264] WLL[263] WLL[262] WLL[261] WLL[260] WLL[259] WLL[258] WLL[257] WLL[256]
+WLL[255] WLL[254] WLL[253] WLL[252] WLL[251] WLL[250] WLL[249] WLL[248] WLL[247] WLL[246]
+WLL[245] WLL[244] WLL[243] WLL[242] WLL[241] WLL[240] WLL[239] WLL[238] WLL[237] WLL[236]
+WLL[235] WLL[234] WLL[233] WLL[232] WLL[231] WLL[230] WLL[229] WLL[228] WLL[227] WLL[226]
+WLL[225] WLL[224] WLL[223] WLL[222] WLL[221] WLL[220] WLL[219] WLL[218] WLL[217] WLL[216]
+WLL[215] WLL[214] WLL[213] WLL[212] WLL[211] WLL[210] WLL[209] WLL[208] WLL[207] WLL[206]
+WLL[205] WLL[204] WLL[203] WLL[202] WLL[201] WLL[200] WLL[199] WLL[198] WLL[197] WLL[196]
+WLL[195] WLL[194] WLL[193] WLL[192] WLL[191] WLL[190] WLL[189] WLL[188] WLL[187] WLL[186]
+WLL[185] WLL[184] WLL[183] WLL[182] WLL[181] WLL[180] WLL[179] WLL[178] WLL[177] WLL[176]
+WLL[175] WLL[174] WLL[173] WLL[172] WLL[171] WLL[170] WLL[169] WLL[168] WLL[167] WLL[166]
+WLL[165] WLL[164] WLL[163] WLL[162] WLL[161] WLL[160] WLL[159] WLL[158] WLL[157] WLL[156]
+WLL[155] WLL[154] WLL[153] WLL[152] WLL[151] WLL[150] WLL[149] WLL[148] WLL[147] WLL[146]
+WLL[145] WLL[144] WLL[143] WLL[142] WLL[141] WLL[140] WLL[139] WLL[138] WLL[137] WLL[136]
+WLL[135] WLL[134] WLL[133] WLL[132] WLL[131] WLL[130] WLL[129] WLL[128] WLL[127] WLL[126]
+WLL[125] WLL[124] WLL[123] WLL[122] WLL[121] WLL[120] WLL[119] WLL[118] WLL[117] WLL[116]
+WLL[115] WLL[114] WLL[113] WLL[112] WLL[111] WLL[110] WLL[109] WLL[108] WLL[107] WLL[106]
+WLL[105] WLL[104] WLL[103] WLL[102] WLL[101] WLL[100] WLL[99] WLL[98] WLL[97] WLL[96]
+WLL[95] WLL[94] WLL[93] WLL[92] WLL[91] WLL[90] WLL[89] WLL[88] WLL[87] WLL[86]
+WLL[85] WLL[84] WLL[83] WLL[82] WLL[81] WLL[80] WLL[79] WLL[78] WLL[77] WLL[76]
+WLL[75] WLL[74] WLL[73] WLL[72] WLL[71] WLL[70] WLL[69] WLL[68] WLL[67] WLL[66]
+WLL[65] WLL[64] WLL[63] WLL[62] WLL[61] WLL[60] WLL[59] WLL[58] WLL[57] WLL[56]
+WLL[55] WLL[54] WLL[53] WLL[52] WLL[51] WLL[50] WLL[49] WLL[48] WLL[47] WLL[46]
+WLL[45] WLL[44] WLL[43] WLL[42] WLL[41] WLL[40] WLL[39] WLL[38] WLL[37] WLL[36]
+WLL[35] WLL[34] WLL[33] WLL[32] WLL[31] WLL[30] WLL[29] WLL[28] WLL[27] WLL[26]
+WLL[25] WLL[24] WLL[23] WLL[22] WLL[21] WLL[20] WLL[19] WLL[18] WLL[17] WLL[16]
+WLL[15] WLL[14] WLL[13] WLL[12] WLL[11] WLL[10] WLL[9] WLL[8] WLL[7] WLL[6]
+WLL[5] WLL[4] WLL[3] WLL[2] WLL[1] WLL[0] YAX YX[7] YX[6] YX[5]
+YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_ARRAY_X512Y16D16_LEFT
XI1 D[31] D[30] D[29] D[28] D[27] D[26] D[25] D[24] D[23] D[22]
+D[21] D[20] D[19] D[18] D[17] D[16] DBL DCTRCLK DCTRCLKX Q[31]
+Q[30] Q[29] Q[28] Q[27] Q[26] Q[25] Q[24] Q[23] Q[22] Q[21]
+Q[20] Q[19] Q[18] Q[17] Q[16] VSS VSS RWLR VSS SACK1
+SACK4 STWL VDD VSS WE WLR[511] WLR[510] WLR[509] WLR[508] WLR[507]
+WLR[506] WLR[505] WLR[504] WLR[503] WLR[502] WLR[501] WLR[500] WLR[499] WLR[498] WLR[497]
+WLR[496] WLR[495] WLR[494] WLR[493] WLR[492] WLR[491] WLR[490] WLR[489] WLR[488] WLR[487]
+WLR[486] WLR[485] WLR[484] WLR[483] WLR[482] WLR[481] WLR[480] WLR[479] WLR[478] WLR[477]
+WLR[476] WLR[475] WLR[474] WLR[473] WLR[472] WLR[471] WLR[470] WLR[469] WLR[468] WLR[467]
+WLR[466] WLR[465] WLR[464] WLR[463] WLR[462] WLR[461] WLR[460] WLR[459] WLR[458] WLR[457]
+WLR[456] WLR[455] WLR[454] WLR[453] WLR[452] WLR[451] WLR[450] WLR[449] WLR[448] WLR[447]
+WLR[446] WLR[445] WLR[444] WLR[443] WLR[442] WLR[441] WLR[440] WLR[439] WLR[438] WLR[437]
+WLR[436] WLR[435] WLR[434] WLR[433] WLR[432] WLR[431] WLR[430] WLR[429] WLR[428] WLR[427]
+WLR[426] WLR[425] WLR[424] WLR[423] WLR[422] WLR[421] WLR[420] WLR[419] WLR[418] WLR[417]
+WLR[416] WLR[415] WLR[414] WLR[413] WLR[412] WLR[411] WLR[410] WLR[409] WLR[408] WLR[407]
+WLR[406] WLR[405] WLR[404] WLR[403] WLR[402] WLR[401] WLR[400] WLR[399] WLR[398] WLR[397]
+WLR[396] WLR[395] WLR[394] WLR[393] WLR[392] WLR[391] WLR[390] WLR[389] WLR[388] WLR[387]
+WLR[386] WLR[385] WLR[384] WLR[383] WLR[382] WLR[381] WLR[380] WLR[379] WLR[378] WLR[377]
+WLR[376] WLR[375] WLR[374] WLR[373] WLR[372] WLR[371] WLR[370] WLR[369] WLR[368] WLR[367]
+WLR[366] WLR[365] WLR[364] WLR[363] WLR[362] WLR[361] WLR[360] WLR[359] WLR[358] WLR[357]
+WLR[356] WLR[355] WLR[354] WLR[353] WLR[352] WLR[351] WLR[350] WLR[349] WLR[348] WLR[347]
+WLR[346] WLR[345] WLR[344] WLR[343] WLR[342] WLR[341] WLR[340] WLR[339] WLR[338] WLR[337]
+WLR[336] WLR[335] WLR[334] WLR[333] WLR[332] WLR[331] WLR[330] WLR[329] WLR[328] WLR[327]
+WLR[326] WLR[325] WLR[324] WLR[323] WLR[322] WLR[321] WLR[320] WLR[319] WLR[318] WLR[317]
+WLR[316] WLR[315] WLR[314] WLR[313] WLR[312] WLR[311] WLR[310] WLR[309] WLR[308] WLR[307]
+WLR[306] WLR[305] WLR[304] WLR[303] WLR[302] WLR[301] WLR[300] WLR[299] WLR[298] WLR[297]
+WLR[296] WLR[295] WLR[294] WLR[293] WLR[292] WLR[291] WLR[290] WLR[289] WLR[288] WLR[287]
+WLR[286] WLR[285] WLR[284] WLR[283] WLR[282] WLR[281] WLR[280] WLR[279] WLR[278] WLR[277]
+WLR[276] WLR[275] WLR[274] WLR[273] WLR[272] WLR[271] WLR[270] WLR[269] WLR[268] WLR[267]
+WLR[266] WLR[265] WLR[264] WLR[263] WLR[262] WLR[261] WLR[260] WLR[259] WLR[258] WLR[257]
+WLR[256] WLR[255] WLR[254] WLR[253] WLR[252] WLR[251] WLR[250] WLR[249] WLR[248] WLR[247]
+WLR[246] WLR[245] WLR[244] WLR[243] WLR[242] WLR[241] WLR[240] WLR[239] WLR[238] WLR[237]
+WLR[236] WLR[235] WLR[234] WLR[233] WLR[232] WLR[231] WLR[230] WLR[229] WLR[228] WLR[227]
+WLR[226] WLR[225] WLR[224] WLR[223] WLR[222] WLR[221] WLR[220] WLR[219] WLR[218] WLR[217]
+WLR[216] WLR[215] WLR[214] WLR[213] WLR[212] WLR[211] WLR[210] WLR[209] WLR[208] WLR[207]
+WLR[206] WLR[205] WLR[204] WLR[203] WLR[202] WLR[201] WLR[200] WLR[199] WLR[198] WLR[197]
+WLR[196] WLR[195] WLR[194] WLR[193] WLR[192] WLR[191] WLR[190] WLR[189] WLR[188] WLR[187]
+WLR[186] WLR[185] WLR[184] WLR[183] WLR[182] WLR[181] WLR[180] WLR[179] WLR[178] WLR[177]
+WLR[176] WLR[175] WLR[174] WLR[173] WLR[172] WLR[171] WLR[170] WLR[169] WLR[168] WLR[167]
+WLR[166] WLR[165] WLR[164] WLR[163] WLR[162] WLR[161] WLR[160] WLR[159] WLR[158] WLR[157]
+WLR[156] WLR[155] WLR[154] WLR[153] WLR[152] WLR[151] WLR[150] WLR[149] WLR[148] WLR[147]
+WLR[146] WLR[145] WLR[144] WLR[143] WLR[142] WLR[141] WLR[140] WLR[139] WLR[138] WLR[137]
+WLR[136] WLR[135] WLR[134] WLR[133] WLR[132] WLR[131] WLR[130] WLR[129] WLR[128] WLR[127]
+WLR[126] WLR[125] WLR[124] WLR[123] WLR[122] WLR[121] WLR[120] WLR[119] WLR[118] WLR[117]
+WLR[116] WLR[115] WLR[114] WLR[113] WLR[112] WLR[111] WLR[110] WLR[109] WLR[108] WLR[107]
+WLR[106] WLR[105] WLR[104] WLR[103] WLR[102] WLR[101] WLR[100] WLR[99] WLR[98] WLR[97]
+WLR[96] WLR[95] WLR[94] WLR[93] WLR[92] WLR[91] WLR[90] WLR[89] WLR[88] WLR[87]
+WLR[86] WLR[85] WLR[84] WLR[83] WLR[82] WLR[81] WLR[80] WLR[79] WLR[78] WLR[77]
+WLR[76] WLR[75] WLR[74] WLR[73] WLR[72] WLR[71] WLR[70] WLR[69] WLR[68] WLR[67]
+WLR[66] WLR[65] WLR[64] WLR[63] WLR[62] WLR[61] WLR[60] WLR[59] WLR[58] WLR[57]
+WLR[56] WLR[55] WLR[54] WLR[53] WLR[52] WLR[51] WLR[50] WLR[49] WLR[48] WLR[47]
+WLR[46] WLR[45] WLR[44] WLR[43] WLR[42] WLR[41] WLR[40] WLR[39] WLR[38] WLR[37]
+WLR[36] WLR[35] WLR[34] WLR[33] WLR[32] WLR[31] WLR[30] WLR[29] WLR[28] WLR[27]
+WLR[26] WLR[25] WLR[24] WLR[23] WLR[22] WLR[21] WLR[20] WLR[19] WLR[18] WLR[17]
+WLR[16] WLR[15] WLR[14] WLR[13] WLR[12] WLR[11] WLR[10] WLR[9] WLR[8] WLR[7]
+WLR[6] WLR[5] WLR[4] WLR[3] WLR[2] WLR[1] WLR[0] YAX YX[7] YX[6]
+YX[5] YX[4] YX[3] YX[2] YX[1] YX[0] ZAS ZASX S55NLLGSPH_X512Y16D32_ARRAY_X512Y16D16_RIGHT
XI2 TIE_LOW VSS VDD S55NLLGSPH_X512Y16D32_TIE_LOW_S
XI3 TIE_HIGH VSS VDD S55NLLGSPH_X512Y16D32_TIE_HIGH_S
XI4 DBL STWL TIE_LOW TIE_HIGH VDD VSS S55NLLGSPH_X512Y16D32_SOP_S
XI5 ACTRCLK ACTRCLKX CEN CLK DCTRCLK DCTRCLKX EMCLK DBL FCKX[7] FCKX[6]
+FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXA[2] PXA[1] PXA[0]
+TIELOW_RDE RWLL RWLR TIE_HIGH TIE_LOW SACK1 SACK4 VDD VSS WE
+WEN A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0]
+YAX YX[7] YX[6] YX[5] YX[4] YX[3] YX[2] YX[1] YX[0] ZAS
+ZASX S55NLLGSPH_X512Y16D32_LOGIC_BASEY16
XI6 A[12] A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3]
+A[2] A[1] A[0] CEN CLK TIELOW_RDE TIE_HIGH TIE_LOW VDD VSS
+WEN S55NLLGSPH_X512Y16D32_S65NLLHSDPH_ESDA12
XI7 VDD VSS TIELOW_RDE S55NLLGSPH_X512Y16D32_TIE_LOW_X2
XI8 EMCLK STWL VDD VSS S55NLLGSPH_X512Y16D32_STWL_DEC
XI9 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXA[1]
+PXB[3] PXB[2] PXB[1] PXB[0] PXC[3] PXC[2] PXC[1] PXC[0] VDD VSS
+WLL[511] WLL[510] WLL[509] WLL[508] WLL[507] WLL[506] WLL[505] WLL[504] WLL[503] WLL[502]
+WLL[501] WLL[500] WLL[499] WLL[498] WLL[497] WLL[496] WLL[495] WLL[494] WLL[493] WLL[492]
+WLL[491] WLL[490] WLL[489] WLL[488] WLL[487] WLL[486] WLL[485] WLL[484] WLL[483] WLL[482]
+WLL[481] WLL[480] WLL[479] WLL[478] WLL[477] WLL[476] WLL[475] WLL[474] WLL[473] WLL[472]
+WLL[471] WLL[470] WLL[469] WLL[468] WLL[467] WLL[466] WLL[465] WLL[464] WLL[463] WLL[462]
+WLL[461] WLL[460] WLL[459] WLL[458] WLL[457] WLL[456] WLL[455] WLL[454] WLL[453] WLL[452]
+WLL[451] WLL[450] WLL[449] WLL[448] WLL[447] WLL[446] WLL[445] WLL[444] WLL[443] WLL[442]
+WLL[441] WLL[440] WLL[439] WLL[438] WLL[437] WLL[436] WLL[435] WLL[434] WLL[433] WLL[432]
+WLL[431] WLL[430] WLL[429] WLL[428] WLL[427] WLL[426] WLL[425] WLL[424] WLL[423] WLL[422]
+WLL[421] WLL[420] WLL[419] WLL[418] WLL[417] WLL[416] WLL[415] WLL[414] WLL[413] WLL[412]
+WLL[411] WLL[410] WLL[409] WLL[408] WLL[407] WLL[406] WLL[405] WLL[404] WLL[403] WLL[402]
+WLL[401] WLL[400] WLL[399] WLL[398] WLL[397] WLL[396] WLL[395] WLL[394] WLL[393] WLL[392]
+WLL[391] WLL[390] WLL[389] WLL[388] WLL[387] WLL[386] WLL[385] WLL[384] WLL[383] WLL[382]
+WLL[381] WLL[380] WLL[379] WLL[378] WLL[377] WLL[376] WLL[375] WLL[374] WLL[373] WLL[372]
+WLL[371] WLL[370] WLL[369] WLL[368] WLL[367] WLL[366] WLL[365] WLL[364] WLL[363] WLL[362]
+WLL[361] WLL[360] WLL[359] WLL[358] WLL[357] WLL[356] WLL[355] WLL[354] WLL[353] WLL[352]
+WLL[351] WLL[350] WLL[349] WLL[348] WLL[347] WLL[346] WLL[345] WLL[344] WLL[343] WLL[342]
+WLL[341] WLL[340] WLL[339] WLL[338] WLL[337] WLL[336] WLL[335] WLL[334] WLL[333] WLL[332]
+WLL[331] WLL[330] WLL[329] WLL[328] WLL[327] WLL[326] WLL[325] WLL[324] WLL[323] WLL[322]
+WLL[321] WLL[320] WLL[319] WLL[318] WLL[317] WLL[316] WLL[315] WLL[314] WLL[313] WLL[312]
+WLL[311] WLL[310] WLL[309] WLL[308] WLL[307] WLL[306] WLL[305] WLL[304] WLL[303] WLL[302]
+WLL[301] WLL[300] WLL[299] WLL[298] WLL[297] WLL[296] WLL[295] WLL[294] WLL[293] WLL[292]
+WLL[291] WLL[290] WLL[289] WLL[288] WLL[287] WLL[286] WLL[285] WLL[284] WLL[283] WLL[282]
+WLL[281] WLL[280] WLL[279] WLL[278] WLL[277] WLL[276] WLL[275] WLL[274] WLL[273] WLL[272]
+WLL[271] WLL[270] WLL[269] WLL[268] WLL[267] WLL[266] WLL[265] WLL[264] WLL[263] WLL[262]
+WLL[261] WLL[260] WLL[259] WLL[258] WLL[257] WLL[256] WLR[511] WLR[510] WLR[509] WLR[508]
+WLR[507] WLR[506] WLR[505] WLR[504] WLR[503] WLR[502] WLR[501] WLR[500] WLR[499] WLR[498]
+WLR[497] WLR[496] WLR[495] WLR[494] WLR[493] WLR[492] WLR[491] WLR[490] WLR[489] WLR[488]
+WLR[487] WLR[486] WLR[485] WLR[484] WLR[483] WLR[482] WLR[481] WLR[480] WLR[479] WLR[478]
+WLR[477] WLR[476] WLR[475] WLR[474] WLR[473] WLR[472] WLR[471] WLR[470] WLR[469] WLR[468]
+WLR[467] WLR[466] WLR[465] WLR[464] WLR[463] WLR[462] WLR[461] WLR[460] WLR[459] WLR[458]
+WLR[457] WLR[456] WLR[455] WLR[454] WLR[453] WLR[452] WLR[451] WLR[450] WLR[449] WLR[448]
+WLR[447] WLR[446] WLR[445] WLR[444] WLR[443] WLR[442] WLR[441] WLR[440] WLR[439] WLR[438]
+WLR[437] WLR[436] WLR[435] WLR[434] WLR[433] WLR[432] WLR[431] WLR[430] WLR[429] WLR[428]
+WLR[427] WLR[426] WLR[425] WLR[424] WLR[423] WLR[422] WLR[421] WLR[420] WLR[419] WLR[418]
+WLR[417] WLR[416] WLR[415] WLR[414] WLR[413] WLR[412] WLR[411] WLR[410] WLR[409] WLR[408]
+WLR[407] WLR[406] WLR[405] WLR[404] WLR[403] WLR[402] WLR[401] WLR[400] WLR[399] WLR[398]
+WLR[397] WLR[396] WLR[395] WLR[394] WLR[393] WLR[392] WLR[391] WLR[390] WLR[389] WLR[388]
+WLR[387] WLR[386] WLR[385] WLR[384] WLR[383] WLR[382] WLR[381] WLR[380] WLR[379] WLR[378]
+WLR[377] WLR[376] WLR[375] WLR[374] WLR[373] WLR[372] WLR[371] WLR[370] WLR[369] WLR[368]
+WLR[367] WLR[366] WLR[365] WLR[364] WLR[363] WLR[362] WLR[361] WLR[360] WLR[359] WLR[358]
+WLR[357] WLR[356] WLR[355] WLR[354] WLR[353] WLR[352] WLR[351] WLR[350] WLR[349] WLR[348]
+WLR[347] WLR[346] WLR[345] WLR[344] WLR[343] WLR[342] WLR[341] WLR[340] WLR[339] WLR[338]
+WLR[337] WLR[336] WLR[335] WLR[334] WLR[333] WLR[332] WLR[331] WLR[330] WLR[329] WLR[328]
+WLR[327] WLR[326] WLR[325] WLR[324] WLR[323] WLR[322] WLR[321] WLR[320] WLR[319] WLR[318]
+WLR[317] WLR[316] WLR[315] WLR[314] WLR[313] WLR[312] WLR[311] WLR[310] WLR[309] WLR[308]
+WLR[307] WLR[306] WLR[305] WLR[304] WLR[303] WLR[302] WLR[301] WLR[300] WLR[299] WLR[298]
+WLR[297] WLR[296] WLR[295] WLR[294] WLR[293] WLR[292] WLR[291] WLR[290] WLR[289] WLR[288]
+WLR[287] WLR[286] WLR[285] WLR[284] WLR[283] WLR[282] WLR[281] WLR[280] WLR[279] WLR[278]
+WLR[277] WLR[276] WLR[275] WLR[274] WLR[273] WLR[272] WLR[271] WLR[270] WLR[269] WLR[268]
+WLR[267] WLR[266] WLR[265] WLR[264] WLR[263] WLR[262] WLR[261] WLR[260] WLR[259] WLR[258]
+WLR[257] WLR[256] S55NLLGSPH_X512Y16D32_XDEC32
XI10 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXA[0]
+PXB[3] PXB[2] PXB[1] PXB[0] PXC[3] PXC[2] PXC[1] PXC[0] VDD VSS
+WLL[255] WLL[254] WLL[253] WLL[252] WLL[251] WLL[250] WLL[249] WLL[248] WLL[247] WLL[246]
+WLL[245] WLL[244] WLL[243] WLL[242] WLL[241] WLL[240] WLL[239] WLL[238] WLL[237] WLL[236]
+WLL[235] WLL[234] WLL[233] WLL[232] WLL[231] WLL[230] WLL[229] WLL[228] WLL[227] WLL[226]
+WLL[225] WLL[224] WLL[223] WLL[222] WLL[221] WLL[220] WLL[219] WLL[218] WLL[217] WLL[216]
+WLL[215] WLL[214] WLL[213] WLL[212] WLL[211] WLL[210] WLL[209] WLL[208] WLL[207] WLL[206]
+WLL[205] WLL[204] WLL[203] WLL[202] WLL[201] WLL[200] WLL[199] WLL[198] WLL[197] WLL[196]
+WLL[195] WLL[194] WLL[193] WLL[192] WLL[191] WLL[190] WLL[189] WLL[188] WLL[187] WLL[186]
+WLL[185] WLL[184] WLL[183] WLL[182] WLL[181] WLL[180] WLL[179] WLL[178] WLL[177] WLL[176]
+WLL[175] WLL[174] WLL[173] WLL[172] WLL[171] WLL[170] WLL[169] WLL[168] WLL[167] WLL[166]
+WLL[165] WLL[164] WLL[163] WLL[162] WLL[161] WLL[160] WLL[159] WLL[158] WLL[157] WLL[156]
+WLL[155] WLL[154] WLL[153] WLL[152] WLL[151] WLL[150] WLL[149] WLL[148] WLL[147] WLL[146]
+WLL[145] WLL[144] WLL[143] WLL[142] WLL[141] WLL[140] WLL[139] WLL[138] WLL[137] WLL[136]
+WLL[135] WLL[134] WLL[133] WLL[132] WLL[131] WLL[130] WLL[129] WLL[128] WLL[127] WLL[126]
+WLL[125] WLL[124] WLL[123] WLL[122] WLL[121] WLL[120] WLL[119] WLL[118] WLL[117] WLL[116]
+WLL[115] WLL[114] WLL[113] WLL[112] WLL[111] WLL[110] WLL[109] WLL[108] WLL[107] WLL[106]
+WLL[105] WLL[104] WLL[103] WLL[102] WLL[101] WLL[100] WLL[99] WLL[98] WLL[97] WLL[96]
+WLL[95] WLL[94] WLL[93] WLL[92] WLL[91] WLL[90] WLL[89] WLL[88] WLL[87] WLL[86]
+WLL[85] WLL[84] WLL[83] WLL[82] WLL[81] WLL[80] WLL[79] WLL[78] WLL[77] WLL[76]
+WLL[75] WLL[74] WLL[73] WLL[72] WLL[71] WLL[70] WLL[69] WLL[68] WLL[67] WLL[66]
+WLL[65] WLL[64] WLL[63] WLL[62] WLL[61] WLL[60] WLL[59] WLL[58] WLL[57] WLL[56]
+WLL[55] WLL[54] WLL[53] WLL[52] WLL[51] WLL[50] WLL[49] WLL[48] WLL[47] WLL[46]
+WLL[45] WLL[44] WLL[43] WLL[42] WLL[41] WLL[40] WLL[39] WLL[38] WLL[37] WLL[36]
+WLL[35] WLL[34] WLL[33] WLL[32] WLL[31] WLL[30] WLL[29] WLL[28] WLL[27] WLL[26]
+WLL[25] WLL[24] WLL[23] WLL[22] WLL[21] WLL[20] WLL[19] WLL[18] WLL[17] WLL[16]
+WLL[15] WLL[14] WLL[13] WLL[12] WLL[11] WLL[10] WLL[9] WLL[8] WLL[7] WLL[6]
+WLL[5] WLL[4] WLL[3] WLL[2] WLL[1] WLL[0] WLR[255] WLR[254] WLR[253] WLR[252]
+WLR[251] WLR[250] WLR[249] WLR[248] WLR[247] WLR[246] WLR[245] WLR[244] WLR[243] WLR[242]
+WLR[241] WLR[240] WLR[239] WLR[238] WLR[237] WLR[236] WLR[235] WLR[234] WLR[233] WLR[232]
+WLR[231] WLR[230] WLR[229] WLR[228] WLR[227] WLR[226] WLR[225] WLR[224] WLR[223] WLR[222]
+WLR[221] WLR[220] WLR[219] WLR[218] WLR[217] WLR[216] WLR[215] WLR[214] WLR[213] WLR[212]
+WLR[211] WLR[210] WLR[209] WLR[208] WLR[207] WLR[206] WLR[205] WLR[204] WLR[203] WLR[202]
+WLR[201] WLR[200] WLR[199] WLR[198] WLR[197] WLR[196] WLR[195] WLR[194] WLR[193] WLR[192]
+WLR[191] WLR[190] WLR[189] WLR[188] WLR[187] WLR[186] WLR[185] WLR[184] WLR[183] WLR[182]
+WLR[181] WLR[180] WLR[179] WLR[178] WLR[177] WLR[176] WLR[175] WLR[174] WLR[173] WLR[172]
+WLR[171] WLR[170] WLR[169] WLR[168] WLR[167] WLR[166] WLR[165] WLR[164] WLR[163] WLR[162]
+WLR[161] WLR[160] WLR[159] WLR[158] WLR[157] WLR[156] WLR[155] WLR[154] WLR[153] WLR[152]
+WLR[151] WLR[150] WLR[149] WLR[148] WLR[147] WLR[146] WLR[145] WLR[144] WLR[143] WLR[142]
+WLR[141] WLR[140] WLR[139] WLR[138] WLR[137] WLR[136] WLR[135] WLR[134] WLR[133] WLR[132]
+WLR[131] WLR[130] WLR[129] WLR[128] WLR[127] WLR[126] WLR[125] WLR[124] WLR[123] WLR[122]
+WLR[121] WLR[120] WLR[119] WLR[118] WLR[117] WLR[116] WLR[115] WLR[114] WLR[113] WLR[112]
+WLR[111] WLR[110] WLR[109] WLR[108] WLR[107] WLR[106] WLR[105] WLR[104] WLR[103] WLR[102]
+WLR[101] WLR[100] WLR[99] WLR[98] WLR[97] WLR[96] WLR[95] WLR[94] WLR[93] WLR[92]
+WLR[91] WLR[90] WLR[89] WLR[88] WLR[87] WLR[86] WLR[85] WLR[84] WLR[83] WLR[82]
+WLR[81] WLR[80] WLR[79] WLR[78] WLR[77] WLR[76] WLR[75] WLR[74] WLR[73] WLR[72]
+WLR[71] WLR[70] WLR[69] WLR[68] WLR[67] WLR[66] WLR[65] WLR[64] WLR[63] WLR[62]
+WLR[61] WLR[60] WLR[59] WLR[58] WLR[57] WLR[56] WLR[55] WLR[54] WLR[53] WLR[52]
+WLR[51] WLR[50] WLR[49] WLR[48] WLR[47] WLR[46] WLR[45] WLR[44] WLR[43] WLR[42]
+WLR[41] WLR[40] WLR[39] WLR[38] WLR[37] WLR[36] WLR[35] WLR[34] WLR[33] WLR[32]
+WLR[31] WLR[30] WLR[29] WLR[28] WLR[27] WLR[26] WLR[25] WLR[24] WLR[23] WLR[22]
+WLR[21] WLR[20] WLR[19] WLR[18] WLR[17] WLR[16] WLR[15] WLR[14] WLR[13] WLR[12]
+WLR[11] WLR[10] WLR[9] WLR[8] WLR[7] WLR[6] WLR[5] WLR[4] WLR[3] WLR[2]
+WLR[1] WLR[0] S55NLLGSPH_X512Y16D32_XDEC32
XI11 A[9] A[10] ACTRCLK ACTRCLKX PXB[3] PXB[2] PXB[1] PXB[0] VDD VSS S55NLLGSPH_X512Y16D32_PX4
XI12 A[11] A[12] ACTRCLK ACTRCLKX PXC[3] PXC[2] PXC[1] PXC[0] VDD VSS S55NLLGSPH_X512Y16D32_PX4
.ENDS
